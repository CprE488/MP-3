XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ur$���c�����X���Zl@�[���؁&�O�����
�Y醂��������_JAw��&�[�*�)i�r�I�����ÜSW�5��L��xK����AՒu�֗]��o��֕'��:}mޕ_k�.�EU&�ٜ�6�k���[�nՒ�.���K��(�f�*A��>�/3��</"�_�r��l�m��×�}��c&^��E$�aR��TS�@�� ��rR� I�����6H�{�Irw{���%�������v.!l #G<\�ǉ��2�0���9h�oCe�%�<���u���NW%�R�`��gl�%l������|��WyQP�Ǫ���
f�(�p��}$����ʭ�V���3΋"x����~�τC3��g�=��*!��rh���������{�Ҡ�`ýz|=�o&���!)�[{�a�X�����uU�I_�^1rҵ����U�ٽ?R���]����R��XI�T��ʌ�甲�+^�X��+���놔pW��#���GЉ�@Y�F#c\�yo���&��s����}�ة\�����	���A<��3�>��\�]L��d��\8њ�'8|��'��>��0}��Ky�7��&Ji�؂��#E튽��	���)Ӯ���& QA%�Y�������������߼%i���	bYcݰO�|K���}s�Ta(��e�*�L� ���a�������L���~�R<���gSpX>Ϗ:��~����D�1��6���/�jXlxVHYEB    3e93    10b0:C�'N,x�R'Q狁b)c��Vv��)����(	ˁN]b?L�!�~�wi{��U����5�⥶0�wWb�Re�	�[����qzS$t��6�@�Ea��
O��t�̀�u{@w���m'Z ������Ȗ�=Gr�z-z�?��I�]�ћX�.�֕J�z��[��?���k���1����Q9p�-B#���Xg�s�A��'I˻�k2��wfYg����w�uX3#Ԧ�E�r�̌��%����ً,H9�XMM�%�^i�	,[9
	��؉Δ�j+U�0jNnOn@=q���w�aT��g����׎�<(a!rq5��
�4Nf5mg�'��.K	C��Y��maI����)�/	�u?nnK�m)�@A��k�mLP��#g���q$\- )�Js�;�>n�m�
���%x��i�K���0�wm� ���X2�i	}a�;�it��W�rJK�.�+т�)[�۶������|�[�u��bf����6�Y6�ӆ��n��B���l�8�7M��5-T��}��]�QWr�i3ZsV��8�CN\��>����s�r��;{�j��k"��X`��wf-�?�[��:D�\�����iU��Ŗ�մы�l�a��������4�I�vg��K��-�%Y�;�y�c��Nt��h֘�F}��93B���C]�ڣ���L�nȩa����F���"�<e�r��r�GL����U��F{|�-���N�Z�3ہA�,=����C��D��0�����G�f��ZlIo��0�%�Y��Sb�bӷs�'IT�>���[���FDOd8�ߠ�_+>b�J�;�_A�6�/'�������8�E���9G�����r���_u�Y�v���oŀ�Z3$�m��jj�s`�b�K��k�����5�K;��x�v{O���*`O����Ő(2�FݶH�W�t"��1?���*V@K��_@L��l 1�*��@2�qhsl�yV�_�{���qQ�hqfd��Wq7j6�G �-xʗ�QT4��+H���w��j�v���Ye����WIx'�}���и�ߟ��H5ad� f�-+³+<��_
�x���rb�aV�#�l�q�!�=�Vzy�=�KW1K Z��(w��]�J�e�R
�6�̌qh�~S�x���G�BC��W
���xO���=�1Ah�`ʍ��4�T�w+)��[��48h�\�|�	����7(Na���7 9�~OG;�'�ب?�SK�4�Z��fO7��qdr�o.:n_6���A!�Y5,���~����i�����煘!����g�s�\h�5�l�>; ��\�,�O�?�k3J���vV#��SueR�#��kv�5�7���0��O����B�GN�\	�J*{¼ϖu Q����g�з�.i[�ܥgC}3���Y�[ܡ��4-/z����L�
�KK�\����&cW�AR��[}ؼ�C����9�}�S�>����l�f��t���yS��՝��?�׏��zq��m�QP!�����l�>�N���Q���(){�D��?v�˶��Ժ�Z�c�*D����<uj�b�0������Q����	H$n1'9�;M��x�Ju*�n����یJrٳ]9��,�@��9��}*�F��ǰ�H�}�I�;�I��6%Uܸ �Z������>wE�&�Ry����}���w�����T�?�Q���4�7����� �G3NەL�r����e�2�oT*��4��y3g��4T�oc5zqL8V�	y����� Oc�%�+�e��A@��k]��e��;+��]����԰�N�8���9���U���;��b���q9v�S�|���]K�VW���r]�S(��*�Y�!�a����8�'��+�~n7^�j�9�J��R��0��@'�Լ��84�T�_A�*C��&����23[��K��^碹����ݨ_Mvp�#K�{-�3� �@�i=�nȑ�bGX5�˫��ղUG����(I�<�t�R+˥a�.�(��;E��!�? @��Ū�j�QA4��fd�	�0��D���J���9����y��Tv���v�&�~"������¬8C�oV�qD��,�p ��m{�$�d�:G�*��_F�*6Z�&^Nٺ�{�`�x"�_�P��ƄB4Co���/�U�Vg*�|�/.(|�I��\���e��j��:��?S�6H�����q���$��ut_\s��/`&���l�1'.28�T�u
�**F�(ۺݘ'�R�T?ꚆN5��-m��	���o��W���gx��}�i6�{⌚��؋���[).��t�\	y	���҅\���0�]:�aK>�F)�S�N�\E,9:�i@5�x��e)��m�@�M>��ٍy����U�S�^;�[~./���F?mY5��cᤱ���K'�x���i!�>���%�8ٕ�% _�*<��3��:�=t��n�s��)sx�tG��*Qb�[�{�n�Ά�q��A	^��$��1[x~�k��->
M�(w��q������c&���>�d�M���}��^�d�^�����C�Ѐ2/�*��u?��C���jՊr#r�YT�8�)3H��N���

A��G�d�[)�|!��A��OV\�V�.��N�֒F����r��U-��૿�	����&�� �U�2W���<�m��KCjw$��ŻXn�����S�|��
G���si�FO^�etf���њ"�v���>!�����_g�fٕ��F�ژ�%���M��<�K��6�QT���Qи��{3��+���w���I�
j�D�	d%���噎�н��e(]Ȕ=�$]K�_���<���`Z(��<O���T�Ŧ�����;�PT���4��AI5����U���)�(�J�5E���;�z:��p���`���V ���#c1ںy���"7�kj�i��u��?5	��+�^2�;:'��v������˲�E��jʦ�<��BJ��L�ri}l"�w"~��`�'=��(�|!�9L�:<�T\�Ʉ�E���1����;J���c�>n(�{��!+����1X��VM��Sf_�Ґ;�`���9a�N� �JL��TK���̈{��ii*��b�ÿI���?[�'���8L\T+؄��~��=n�:�`���5L�{�t�;��5RMC�"��X�L����_�^UG�O���]��p�b�{�#�oe9r,}z�$�p�U���ꈡ^�^�	�;�pG9�څ��}���|�[K9�V�\��3 ��=@������S��>�Y�z���j��.>aR��� �9x�yS���Zxr��J�Uc}�Aa�M�)LH�� ��ʳ���"iED	bI����WNb>��_�vF�IU�Gy찪>����8:�PȊy�=�0�����C���!��,�0V#���.HrV��A�*ކf�q1�2
�pl�7��+褚Y������`R��b�`��[�Hس?��Z92H���-=O9��h:fB;���'��7B�d���^/��d?ؓ��[�>��*������[��u�:(z���	q�5��A<V%�'O��)a��3n��p�+l�8t�.���w��0���8������"���3�Sk���,Yy�1�ľ��֛<_/���?�C�e�fұ�ӼĬ{����>bd@�!$��EU�Y&|��)�m�!�"�s�R�j������ %E�gtZS������`~�ޮ���_�:��Z�rC��>`�H��M�(��mT�ՙ}�
�)s�+'�FA��E[q�L�9J��5[k7ir�&���'�;���&9T�!_|&���o�=M�t�|��� c�z�.��`��[�**��]�>���p`�u1���	C��0����%���h[���Z3ö"F*�T�=�w��g��W��G�Zͤ����T���<�,���<V�N��{?���(��~ ������ �=f������h��,O7����iJ�O�iĺ��$�Ke#Ӏe�X�vmhL�=�R3�l�jM�9��}`J=�j]wy!�qHcQ��;�C����B-jИ@�{j�V�����qM:�r'��HxZ���1��q�{ʑ�T�[z�v5͠���*ދ�v$���2EZ�
�:��>�yC������ɸ��݉�!xH�R}V��
Fyi A�=�_�U2WN��.@��O��C.t����c�