XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���X�Vܭ1� ����T��52�%@zt�,"v��8�����|���}h��?��X΄��q`U��-D�CrD����#c+_��ײ�+r��	�u���x����߰`/�u|Of�TB^6� ��Mޭ��.E؄��R�Fs-�ah�.��喬��(�IY?�yV$x��7L�=I����%}k��\>�D�T5��_�+��(x��Ћ>�
C+�[++�~��´K�`|v�\ʧ�ص ���`'�x��:+b�=�;!!�����ԎD��r�͹%�҂��X���(�:��L�fT�jQ��!e���a;�F�=,�m팱�(J�aG"Yy��r,�!ҡ���{(	z�UH4m�����Y�֢����Q���6�T=���a�̳�\g�KK�@�`��\�� z�Ĵ�
#��׈�:�ç۹�.$�M���#r����U��e�N3_I�d�
�5^���1��@.,��MD>��96#ܧ(�� #�:�����%5oh�K�4픦]�' �>��#`�������g҆�U��ͱ�|�	y� _[�g$;�Q>��V&�()�p��x��N�c5G\-~o����Ba��R$���ϭL��`�������@K>��&z�����ddc �o�7��vD���9�y.�}���j�i`��Txȇ:B2g�[N)��֠���܋7H��2w��� م߆���ݧ-S�M�pwP �]A+zЯ�9�]�U��;-B��(�-AW��so��k�wg�XlxVHYEB    da59    2e30��hT�?�֨�	Y���.<�[Re�*� ��1.�Q�0�Y/\����r�eH������i/ļm_��	��G��hyKn0O4�^��)�飸��,�	a�<�Y|ڏG��(�{J��� ����Oܠ/M�	�c�E�(�u��_�KC?�LVJ�y��MW`��=����s|ӏ�]&���]0�ږ���4f�0�im-�V������P��p8����]q0P`3�Y"1�u��BM��u��#��6�y���w�L~@<�~����A8?��/\1+��#F?@���|f΂�C��/ 10s�ެ3�9�5־�K��3��lך!�ۡ�LXeK'�5�z(.vC{�sZF	[�K;g�s.&8�k��a]�-D�M�X����p�ޅ.X
/��w�^4!�7,~
�R���8j��r���SܑM�q�r���r$uZ}n�D���������O!H�h/��9��� >e���:�a �!����Ҕ�y/##�H���k��i�na��=ŢRd��o݋W�5$�f�D�\N2<X�MD8��);�e�E��E=��S,j5�T�O:ݹ[�Oۇ&ϵ��6�cNP�<��7{��|-g�W����i�ۤ���5뚩�����6{�DFpz�zX���ʨ)�,ۘ3�}�/���s�M�Mz#��[�/j,Cm�Rw=���e��X�I|�i�C<0�/�V�ɋ*>w�wO`:l<<gi*�8�P��2�!�Y��f4�@sVB�1�=�y�#�����m�֣�՘o)!�H��dF�(����Jk+uB�����zܨɍ��mEMY���b!����&�x9��$r%ӌ^�g���yoR�K���.Κ�����Nvިv	L��	ݾ�r$�n��o�-�*o��h�xt�����~��Y� wt���h��7O�9��z�}tߞVZP4�9op�3G��Q���Ѯ.���S�ǻ�S�L��ؒ���7��:L��K�3�3�I/K���Z��Y�<:�����w�H�'66G�������ƪ�1U������Y0�S���֫r,Ӯ$��l�v�T����.�s�jI�����9I����f�	m�^A����=!y,8���˖�6j�r{��@7�\w}��]������R�o%F�C���ؓ�	|��;V��'��+�?LC췽"�E� ��@�\m��9W:	��`��rO�?�����35�E� �j�ۂ��������Uf� >Bo���P���}}|�@@�Z�c�� ����Kx��T5`=u��B�y�eWp:�|2�����Ɯ�q8_���.�2�Eq����?'Z<
�Y�F�m�(mÞ�����U$6TI��ɐ���4c���D��'�Ï�Hl[/��z W�W�@�8�p:�B�@��D�\C�e$:Ԧ��pR��8�j��LC����y��6��!�d�x�7}i��q��|����}�Z�HOU#�S����WH76�dv����� �-������#[��sQY0Q�(��.�e8ג~���[y����6V�{�74�ie��F���YP>��~>?�m"ծ��xr]h��-d��C�3���9�ptY�^of0��<7���������A�r*�-O�Sŵ��	*?�J������Ӏ��P�#����	:��"�O0�|�j+3A	00[��YLn�ɛ�YL|2��LA7�=8W��a�S��d�/�\>���,g����e~�F+��Yu��!����2��"u��S����8����c���tj-����|�C߂o�B�@�SIg��\�8�ɢ��7�E��p�d������z�� ��]j�u	r��=QH�3h��$�[�/{�A<�)�����y�zY��\[j����qpu�S��Q(��xjʙ�7�M�O/},f��nO�����ٽ���W�8��I��_+�m���~�
���r���p�֘�y�W6��,
��������$�omٶ/>g��NRy��<}���X�R(D�q[<��tJA�{����ecC�F�}l��6��Ʌ���q�(A�e��C���P�`�����0��S$T��:�j�l��W�~�gVf��mR,�.� �1)�[���Q�^�n�]LMê��&>_?:!t����8Iτ4���/���>�+����<v�]%25�����gF��	��/�n�c�&�gV�;�ޖ�����\[k.4z�Zǩ2J8�Ü���tƖfY�K"�Z���C �/4�Ja){Z��q(U��[�Jv*	�sk����x?��f�wZ��#K�NK$g#�K����F|kB�?�fֆ++ U�bz����[�Y�/�Ѕg��O�X�]����<M��HH��G����u09d�x�y��vv�N�����#��+Q\�ph��s���g��N�g8M2�`�U1UP#(c~D�V�g��.�ce���Oޖp)_��H�+Q��<ӣ��?+Yca�=B�G�~h���3i�ic�,�D��ԒjT��(���qOq�<&�v���?��m�G��9�]���B%�<i~������뎎���[�/�F���8�zւ���#^1�e`��}_�K�r2c#�̼d�6[��3�9(Ad1BC�wϨġi�5�����|�+��P�>��h��l��֊���U��"M����^TVZ�����N���M��]�Qq].p��QtN�F|�����	-U��R��p��A���gx������悔�6�Ί�L(�>v%��&ļ���$�`�Q��a6a�7/؆v�Aݫ8��r� {l4@.^MQ��V�n���x!wK�w�&k�s��bo��"n�_1Vy8]��$��l��Rh�K��b��Е�g%����U�۸���?և�%�S�C#4�g�D��%d��r�����h��t������^v�Xmò�,h�l�b�~�M�ZB���I�z�>���Jks�a�(�"b�['r__maA��@�C˂�k2;�l�(^�8�����"���7)�[E:��R;cr�`AC�Db�Y��6O���kM�\�c��q$c����ַ��Q�"�ps��Z��¿l��hRl�``�"Y'+�sZ2ԍ�|�|��{��HtN���O���e#��-��t���m���(A�Ԩ����g*�cDu��^�LV���9[�����c�o�59 -@ļ�� I�����41��/��@0�E�����������V3����tu/���/���:%��/G���}j��B�w��¹��@7�K��W�0D����Qp�7�S��=Ԝ�'[Vw��'������8��	+5 `=a3U:�����=�`�[5�xN^�ͳ�EH��c>x wL��������i%�J=�kFW��Ui��>�����-��u��*����$�%��p�	D�����W;)�+�]I��5��M�����E��q�k����VHu��9�)����Np�+E�޲���&�.�L��H:�7�q�S_�I�N-0��+2t�T�����=��D���0�ø֩`2�>+��b1��Bw�t.	�	w���圌ڞ��	y�w�ȳ����1d;_Ըn��$7/{�OV[���)DD)ӹ��LGFK1���??��2����^�HT�W��a�S�2"�`�\�~E���u|S�� �8�K���Q)�>���1�xK�-VX�$��)mN�6D��"����hB�'�䲤�6;�LZ>(M�xWYg���ܹ��(��nX�K�®��K^?�qQo{ԑ�.�f�����$�g��u܋�2�E�~��5�j��8p��!�M��k����l�(�!�S���u�r#�������j�Y6���ot���9�ڜU���G�T��@U�*��e>�(Lc����xѝ,JU~�!��!�#t7G�Y�S����ci�=\X�j:�(�[l`����	�eB��"�E��MÎ�s^N���k��#����c����b��fUm)���Z�g��0/���y�ygw��2Z���H	��\Jw[7��gᲄ�U�'p�։���&����ʱO�P�B�����u)+ y+�F:okǡE]���نK썡i9.kX0���ԩ��֫�����(��&� ����&3־�Ǡ�$��LfV�K4������VQ�UE �t��	LEJѕ)�����i|
�F� vz��bϙ�{	R���^	�#�&�5�>�p�Δ�>Ns|�cdm�3��&Jn4�"���hqn�o����$sBjR�OZWVu���*$i�x�ƴ����qD_5[���M�8����
��)�,�YΛ벡��%�j�ڠ($N>�hms}��m��7��ad�O�������s#p��ٌoo[�������qV����l��Y�e��'�_<�M`���7͡��J\�u�7��a�#x"�WZ�)+��i�1B{�*���5��� ^!rod��^y������!�����fF|>��Yc�UG�ޤ�Y#�|P�*O�DVq���YM����ص�K¹I���V$&�
&��OQ�	���t>WF���%K>ӷn}�d��?2���D�f%�x��a]�A̼(uV}iO�Z}���s�6�3�>�5�Y<>��X!�D�i8J�M��n���M���"�d�Զ�>��A��"�0�62�޻�=���g��Q���fQj�Nm�h?�P|r�3�~�Pٗ�x��)��	���ϊ�_m�>Hw���Q��P-R�[u�I���f8ܞ��0�h� o�^e�"�pptqC�g�/1ؾ捧ش�'�q�f���`�2{$�I���<���(�iq�׸��q%m�&�ϗ�������1u�Qt_`Xʇ,^���!���Z��O1�f>�O�ck�f!��{}��bk8��'��q� ɍ�N��z��YTeR������������6U ���2����!�-%��&@�$H�!��tsވb8��!8���G]�ڱz�����j�>;$0�B>�������А��F��ޅ��G��t-�x�ib�Ӡ���}����S�v5Z�%E�ӳ8��1W|�x_�SS�Q*�Xs3Y���cx��l�tyq �Ղ��>�n3q�G�?4��u_/�,V��L��g�v�E֫��?�PY#f���ê��1GBſ�	�p0�^:hzm�+��R�����?7��1�p�����q�p!�:UZI�pȰ��.�}dǲ¥a����W�$�m�G��͛�J��w�7��Ucv�
�xO��3�1/oи����Yv�3w�g�S�����P�xhB�^�
����g�wx�t>C�yG��Է�xe�^� 8s��W�s�ӧsk����<Rap�z]��?_�P�5;T�m�ZH�n����W|`�^7B���k_+BUo����[��ԋRX>P��e��;.�Q�Q����]�0�����g��E��^�x��)���s$���1��: M�ȋ�>4�w��z��!���[�I�	���3�qt_z�2�"����5r�cX��Ă��Z�Z�@�K�B�/姈��D.�d��ZX*��rW{�-{*t �V(����^�v��[�����1�ԯ�z�8%!�	Z�O/�8�5ԋ�i,�ρ�7�:,Je��N�}�6i�F����O�K����g�-u���*v���=�e�ڇ	ɖ�G�{��A�n:�A�N�D(��IR�:c���~{�B�KS�H r��nۤk�Q|��	��%����j�9]k�WN��N��x��(��_@i1���y��ڏ��{ez�T��Jp��y�.@/��n��"���������5Cj{��~�ֺ�rX�����Y���0���v��aL�v���
��&�!:X�1��Ɗ�(�{t��n�yJ&�.���B�o��YM�9��<�$m�[c���,��z���`���I�4a����*�18l=Xs(ii�(�0�C2p��&^ka�ho����Z�웻�뼁����+����?��lp!�zW�r��=�E��в���� \�E�*<�ހ���o�R�wz�c���'��%'[�R�3Adܗ�3 ��u��aQV
A���~��F�ieg,y��SK������ӂzH��ё�ƈ%N�A�(6U��+�׹eqOk+�b��R��A��i�����:����q�Iw�+��e�8�k����Ɗ�����EQR�8t"��MSn����I�T+%��6� ���Z��g�5�~��t5o"Y�l>����g����V&�H�2�3�(�PN�0�J����B�G�\� �-T��V�9U=��?xR�u)6����G*;��鹓��|Y���qP��r�x�ƺ��[�&ORJhYz 	��߰E�GR���M���>6��02ц����(I("���I+׍�y3���&�s��RGb\���"�দq*��h�忘X��"��}�T����ʱY��j��![�w�5�'ޝ2Z�0�
Ĭ�G�]�;j��40փ4"$�J+��/�퇾?V�A�:A��B������!(��P!I�&�)��F��.�O�G����*а�y�uN�	x����"ǻ��n\�M�&Cu�G��=�{!Q����]���vn�ԓ�qZF-^��Y�i�$r��]W/�fY��� 3�Ή�A�k��'Q8sM��| y[9�![����n
m�O_�5宐�e {�����DG�l�pG&[�q-H�ܥ�T�չ{�w�·��ˇ��g=�0	_������r�����V2��#u�ѧ���눓_s��@��8��P��^mF���y�� �y붘w���h��T�ؕ#6��+���Ŏ0e������3�V��P��GO���A}x��g�B"���a�$��m��D�陭��I�.�����ZB-� �#���̡�Jʉ6a�Ȓe L�"����kU��,��0r���v�y/%�����92��$Ja�|rc<��'�1��#�����^z'Qv�,������(t.l�����)��Z!x!l��-��:�i�TC!E�Wq��v���,ӝ(Tŋ���esf��4��,�(�Џ�du�[
q������1��h/&�B���M�����Yvݭ�r�D���{�=���N�F�o��'��;�27�=�Hu����P>�e�˰b7X�>>6N�kki�������{I�C#�6��^�Ӻ�-�;H�n�e����e2���-q�6�3�EK�_�̖ihc>s�Yʻ��J�����t��(c��3����<�	���/��ܡB�uv�N�����%K��rc�xH�K��Fu�rFh�!�I�*�=x`axY�(�ny|	��"*	4C�����OQ��|da�x������^���'�O�.��]Y^NS��e_���xn��|co-���D�� �=����%���xw�L˿D@Y�pA8�n2o,����M):Oݰ���s���~���(�@��A��b��;q�1UU�JY�+^<�I�{[��'~q���Y�����L�,�c0��3�QE| ��Օ3O]������bR����	����8,�֑z7ɱ�����V����x���:���GLk�{�H���Ļ�d���,g��yA�Z(��g�����>�&u}�Xr'��!��fJ-���$K��ݺ[��RH���J� �(#XN���HL�����PC���\�Oל8gP�P�(b,n.OL��@Z��������ҧX�%�(O�)�Ո�O��sp1��f-yj��?�mhO����"G�0�i��(f�.l^���F��W��혐��*���bg&X�����g�g&���ːt�~
fO*U`��c젍W�mA6 yo�j��V�.3�-N�ڡ�g�����%�c�|�/=#�G�Ƣ�^�(�0Iir.b��B�j���\I�%����f�A�=gc�Cac����B/�Ǩ!���k]qj���%ז��O�	�'��+��3J�I��3���pϥ��hT��ю���Ax9h��D��R>_�rJ�bޢ�%��S�
A��V��Y�M�KMyc�l��k~��PF����yIOU50 @����\�� � ��P ]CQ�U���0D��=Y�Q�k��� ۖk\�;�C�6�u�l���b]>?�̄���h���6�2D5��JA��1xB�@*�Hsq�ǌ���8�?M2��ӆH�v�����_�d��2y�y*E�W
��ؖ��F$L�Ʀ��:������i���������oDNG����!b ��} �bDc$~Է�>�u
{����{��Ty�n��.�w�j��8��&�����8<�g�-��g���N� 1���ە]�Dd���n��������q�����h�u�𑇶��\��:����C��|���[߬B��m*��	`m�������7��ռ��'\��y����tͳ����{�;�<!����<���o�̟ؽ,9�9+�Q�PY��#Nβs�H�hђ��R���<3�ޘq�,��t��=�KA�Oao�v���3ĵ_ԟ#����vjR��ޜJ�j��?#�،(�~|���L|��D��+1f*旯���;�@��s�l����r���\z�Z�F�m��ulN���HM8��AWW�$�}������V�����JhT��\��S����!�PCX���_�f��q�aL�,���0�\��Jy4X?0�3H]D��j�������� A:�A!9ō�-�3mg7j�%h��&�W_fN'3jޝ𿦷�l;�)|�I \#�����m�/��*}"����3su'1?t
�����p�P�?�4"�o`����|�E	����	�4Qa�����i��Cge`G��߼����;f��	�(�-ܞ��R-X����O��j�Fl��] �sE쉸��,�`PF
kx�G3'�h�B't�A��CC���|)��=��Y3�ܕ��R|��<�ćk&��E�ׯN��7�I�ǳE��]���D?��`�M����M��i�Z����4���	���j�QC�N}E�T-��ّo6�Q�lC2$K�p �b<������5���IShG�Q��.���s@�J1����n���	���#��}R���9ﭶ�6-ȣ��$�hlF�SL Q��Q`�OnF�{}��$��������_��1ţ�����*b�g�Y%��e�dQ����EBD0�Tv�Y@�T��}�d� $�Aָ@�a5Ağ\�r}Yl	�<�m
�	�!|�hW�E�u��]�QЁ����� �K�+$��{,��;��h�k��f4(��ז0�g�#�7n����w�C��k�������6Yɐ�D���k1����[=�π^��۾푮�Z���q7���!�i\b�W{2�F׊��&��E�d� &茤a!�Wqj1�M9���>��@s�����)��-[�/������g4H+/՗'h�;���>Ly����Xnd��l*79��&x�Y� ���Y�gi� 0�gQ5�I�q�~�+Ǉ ���(�/6Pu�DC����I��+x*<ɇ����t�pK����f��=�#a���W��7 �^��st�EFs(D����`fr�I|�TA^�3�!�+��(ܧ�j�#Ģ�ł!b̧i�,�Y��V�E|�u�2�>z޼��T7�
"��U+͓ն�S��:�}�]��Q<
f]N�+���?.��v��Xp�F1T�D}	�P���-��4)�~&�<S�/�k���A�r�G��p���gR2lR%�S�OR��}���p�N�ޮPW�+H_��X�1hՐ>�I��������(C�?��0�O���1��un I}jl�O�d�����G�_ǌrn�`j8����_j	���L(2 �A��Fc�����w:[�IA��xqh��FY�M�t���
J�sj}5i5Mp���s�!�3O,�)�2�KF�y	C}Ԥ�2�زF�j����2U)��hU��u(��g��(1�<5:�0�Ȯ��j�g�]��E`}W {�K����G��	��ȧuP���X-����{���P���m�����"�����i�g�K�{�O/y�.��Ge�m�Ç<�Hh"�`E�e��:����Y��g���� R,�ճ���Vv\vO��0έR~0"5�[#�-:�(����m��>�"Ϸ�(�uU�"J�[Cn�$�4�ռ
�@��x����s�ʀ��n�\#���i]|M�äBQl��2-ڊ�:�]jo��2�^O�}�է6	�dˋh8�L؃�Ͷ;җy���4�-��f��m1r�)��硛i�9�b�|�)?M0V�d�Z	�)T��U���a��q�Xڲ&]����r:5�BΖ�.�8щc�[����ǲ�!V�1�؇�:m��%,t`����b�7�c�d��=2�|Tߌ�4�<Ғ���b\Q�\���y��q��
 �(�ڏ���-)]bF�l|d�KV���'��A6JM%A�	 �+"#}����q��
��ݣ5m~���=%�cdRޘ��>�LJ,R�um���Z9�)�^�+����V��'O���p��0w��A��qP���'��aCȗh[%{c�3j��F?�@��A�����KJX;b*�h��D?��_ѵ6JN�-��¯�>A�w�R^M�f���Y\���d��%`O�D~y� �$J�4�\�F'�qo�i�O�h+�	X���Ѽ�7XM!v
���S�N��F ��f&�Y*���W��k�^�`��)$ m�� a���w�ZFR֩R���� R|���n�Y�c/� dI���uJMԌ����Kg�g�Q���y#�AM�Sѽ���\�Bs�aC5ݍH�d���#�}I�i��P�hdw+���g�HuW׵��r`��_���QQ~���m9�������`�I�Bn�MFqIDi\���v&0��Bo�"��}��L*,��q丘$EV7�Ȋ�쓉:����(;~O�'�N�}wޞc:-�MS��S���[��޶���-�﮼1����\wq��/��vk�н�ĭ4���ZO���j�^�U!ѣuִ���Sc~���'J��%�|?����j��EqK,�\
[��nQ��X�� ��@�j���n�ם�{�}�p��y9�c�8�l��c��_W��H���t[�(���T̛�J�eH��O$�t8萘��1o�C�����ld�ً�?"4�u���'�Z�����QrL;F�l]]�N����Ґ���<�������yJ�, :-ڼ����>	OzCJ�&B�>kg���2-8;.��@���v.�܈ofw��G���h�M�엳T�L�E�w�
#�R�ۨ�"1�����I�#���0�}{����E���#�!�ۡ����BNS�/7��W;�����[S�N.q}"��|"C)j�EP�)���^x�����݆�ZI4�[R�I���?�� �={;|C�t�I�G�q�94�@�d��b�$)�9��H�SO�v��Z�7�*�+���uW[��-z��nL�Ɋ0=}�e
,[YE_O]T�Ό�HB4J�V�����R���zM�`) V�jjˀ&K��c�|��$�_ͣ�ԕ�M��^��MV'�-� ���ߒ�5M�ig��=�����_]���E9=%oTi]�(R�i.	�|&j�*� ���Ed��-�ml�bT����JU�