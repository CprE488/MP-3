XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��X��7ލ�N>H/���=���(_�XU��^������z}�]��Q<��:@�{
A2� :u��Lx�\�%Bc��`֎�I6)� �ԉNWVkm:���{������W5�n��=��,�ީ��P,���Kk�0y�0�@��)_�D��I��d��+Z�h�r��5���u� %G%�'d���m���:vD�%���vO`}U}�p;ȋ�k�uf������al{C1�X���XpNŐ|���� �O�e�Q쀸�a���X�IO�ݕ���f|&�����"��$�彨 ��w�N�cm��$f�p���(A[<2���:�rj2�q��Ll,�3���hW�k��
�~���qX��u�.�rv;��ra��.D!�PF�#>�h$.�&�XR�I�t�(4l�6�����v ���r����:�^�����<��_?�Ξ�qԂ����Y�"�� >߄�gӗ?eV��H�|�3�2{z�@Ѣ9�C�6D�TG*�=�,���B	C�ň� |���{3���9�LU
H8ר��8L}T�~�y����gvX�~ȗ8`9������k�X������]#L�Ѱk?�~�f2E��.�R����wo�1%}"r�����УD��'k�XFw��kfό8X�F��7�Y�=�66�b�B�v��iH���.N���A3���",�l�5{&8��%̣	T�؇I< X�����&D��V����A��D�3�JFۢ��_�s��U�Ja߰w0bd%�U4�S�XlxVHYEB    17d8     890K�6|/�?{ ��\R��f,�c���<e�0� ���u�	>�%kM�oq+!x�N@���r�5-��DR�]���q/����m����5�Wb[�π�b�Ym�����	_�X-����T3�J�1ȷ��dAea9H� %�f��_�
�Ȏ�?�ޡ�� e����fE�M���ƞ&��w%Ի������rROֺz�[Ծ����ԎsH��C���_��ɸo���� ��wb��T��*�~����نe|l�.�"�vzɰ�H��ꈕ�Q:Fa����k&� o%���5���s�g�����~��Ғ�{���[�k���n!_E�K2�3���Two~CӃ3u��Ķ� �1K1W�W�v�R��<�W*ޞe�6'�7�E���gaT裙��95bz;�Q^�?����w�@%~�~���ѿ<��:�+i�!���?�DA����7��y���6��}�x* �dZ��`�%+�*����ʣ�EV�u��"����^��A��[��3�H�������`v\�k��h0�n%��dx��v���ɹ�Z����B����A�v#�N`B�Z����J 8-�ڑ�`��^�n}=�F��� m$���O�MX�H�����p�+ԛ*L����E)[�U�X�)�O��?��4����?�/�H��w�4E�4��G����ѻo�7��l9yS�5�7�9 <¹�54��%ɟ���5Y����\I��H�>�զx��i��
=��/�O�:��ٚ�$��nLh�R7��<���Y�j�,Tt�8\t�bѪ�g����v{���&����د�*Bj���It�[�0T��,
�MyEE>������ ��_F��1��*֛XBܑZ�HtGѳ�|jXY���zi�O��Fvn���_��S8E�I~H�Z�b�8wN������������, ?�]�׬oy
vB0fr�g����P
�������;�].���b&b0��Z̨��*���UsG@�wQ�s4Z‘���~2nK�3q��P_G���m�3<YA��"y�4Q���5����~��^�p�,�^)ϑ��Me7�qň2~V{�dw�@cS���"�{����ٿ��J�p��|KIR�41���c�7�7��eI嵋(��dWI�ǳ�SO$w��N���R����)/�-��_}&>�Cc�tq&�c���߰���c���� gG��wE*�A��_ks�NWx>�=��Rc���	<�}B�#rm�G��Bp���$�$�C�7={�3��闚��Y�'V���U d��[R���3{dɵ��n^_W^��l�\;5�,����:�#�y+�wi�'�J�N�$��]h�Ǒ�(UA� �����i�"�5�'CqV1�T5j+W�x%���oE�����X�E������j�-�M� ��" ���˷�w:+�]6(.����Rq._Vn DXJ��X�A4��d�;%:>���|q�$�}�~�Zd��T/�0_�z��f�E��W���D�U���k}'�=���W�<E��ߊ�3�����T��R�"����a��c!\���.���F&�V�H�B2W`ݫq Q�˶��0^�#j����O�0ߎV�[R4��C:��!)o%Y�|z�����-:8���|��ce�6���W7� hr���ĥd�,��+��:&��A��>�B�vS���$C����?�:$L,sS�Z�H
��9lZ`�@h���J���CGV��z�	�=�`w�1�҇,�;�shr���vs͵jm Y�(�3}|l�����d�,>:������|����?�֫.�?Gd�����L��l?eR`�Sn��>��!������H%l��"I��޲J��YӍ�(I�T��� ���i��m�L"�E�$�Ԩ��x�m;>d�O�=�(j�~�x��כc��\c;S�����W6��u�Q�Øɨ�]+z��tuJ��-ٳ���Z ��!��h~�׻����`��[�� c���xUؘ��KE-�,%�<N�M�>-�ъ7v�ۆAjZvl��
SBX�K"E�Ӊ���B��|����+���nh��7�'-{�!���2�yA��u $�F6�t�c�&)�q1�F+�v�����ͦ�����B�g��i����JdHg[X����xɯ]�� `2