XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����?�N��v�Q3|,޴%�J�V�e�8}���G����T�i:��֏IS\����i�.�F��mxy��S|ɐ��SV��#��`@�v��y��$H�<"�La�c�V��$����n6���`j���V�=����=#�i�C�]���%����GԠ�X��u>tR�x�X$̏� ��뚔L D�����/����%�YQG�7~HK����}Ke%����E��Xc3�R�p����	1p��p�"�F��I������ �͇�����o�SM���SE?� ���C���d�q(w�ڊܩ}l�Jkkd���Ci3�c[(r/��5�
�3[��:L��HǊ��Nz�fUF!�}��;�4$��8�с�m?���A7\e�l�Cä@�H4��+�˔��ZAU(���gZ�澬&0�I3�$�w�!�K=��4o��zy�tl͉�/7{��ql{�9N�`�q���)�4��x��gm����e�A&?]}�=?y���k�H�H��x�5!��S��(df�}7*��&qBHZ�Aszt��B�����&�_�gZ�P#�*���|��V�huH�(-��E�#|?0
��sQ?�9���F����|��$ˎ*m��J,��_��C�:Ҷ�R_'����K�>�Q>-B����$L�Qr8�[���!l�b���!��U���|ȦYj��.=:q��9=���X���!bxۿ��9��@n��܇�N� .Bi�c0;S}6{ϼh^� .+	%g�6�!B��XlxVHYEB    15b2     890;+��ٿǌ��Ŋ3����q��V�K��4]R��v��b�A9V_�)����2r�ex�ǓKc��۬�4~y�F<t�i������˜{�V2Ko��	 �r�in�����V�3��MbF+���X&���Y1ƞ�М߫����G��@ys�2�˘3�r�	o�ƃb�f<ΐ��**���L���|l���9p+�[��5ˆh9}������df�k�활�������e�&�v�T���Dr�SFl�_c����f�8� ���ܧ�N���c*�N��� ��</��{� *\wpl���LoƟ3��֔�O���'f���)j���;�
Fg�t�D �A�iӹ��W���iW�P����Ÿ��N����ZYĝ���U��:�M�{ũQ;
'�L������0(@�Ε]pq�����;��e(�q��{�Z�#,�32��lD�߂�p�2	K��!Hm�:t��(��&�����w���R��(|�����f�fx���v2���� R�%�,��=��I�)%��ݳ�ǃ�5��	^�'���6�9t����I�؄i/��S�\(9�hKƺ�-㤫�	�&!����ͩ��y�M'p�
�������	|`���5#��Y�����<�(���p�F����0�� �m"eN�7�S��av�fJ��#z�>�6�>�4��Z��)]�U�Z�1�2LH�]�l#��2����U�d��f��y��i$!��|�+��ِA>ek�%F��zޚ�u�FC�Q����H^n�6�*3�HQk�����B��5�f�3un�Xx�mn���-����7���{��s��M���܋%>�B�1���Ed�_�ȧJ��5���7�m"�<0��ڭ�M��P�&뢋,ڮi��'FuH���/k���~�$e���H���Dnb�pel��)�����>�I:̔����Bߌ�?����S8�����ؑ�頱lu�c��ּ��b�3�l'�)�G-��s�$�H	�d��&s�ma2b��1+�l�r �@l`ǁ��*d/�
n�uvsw����0�8<{k��~�Uj�� �)�_�hX`a�i�<bI�l!p���>4�}�;F�?��O'��yy%��jڏ�~#�Q$X�����O���\)��I퓄Hs3��\}b�	�I�+R�Z��[k�h�>�����W��f�>�Kt���f�_�����t�t�PYo�N���$�w�݋Z�%jHcCa\�d���ۮ'8R�µq��8mUdʄd�����V�r���5�G#�4^:��
���u�����I����/�b��01�7��%�^�yC�v����䶽f�-�ڛj��(G�o0(��34�����z9@"8��hL���0��g�!%w��d'�`0?��#�=�qg�n��(��f�EE���qb�����5B�d��[��v�PG~��tC/���d��a�f�n�_h��WŌMί�鉥#$!Rށc�D����̮{��8��M��n�b9��=��E+ l6g�\8��3 !��'±�U��N�{ܲ�.褛*� ��hS��p�xTa�=]���fҺ�������^>��a���Ƀw�\k�( 7�
N����2�J}����v��=���S!p?��N�Y��c�r�%�ql�!fn��c�7�h,(�-���jǵjY%`�.C=@�5��N-[�-��7�%�a-�#쀲��]a�.�����0�����)�>ߓp��+B������V�mW�j%�~S�S8�Ɋ��`��ځ�Y������(w����\Ħݰ��U�R�W�7`4O��+�G���v�1}��N
��J�R�����`^O>a�����Fd�W/E!���.]��;��NC�[�1�y:Y4d���k�&�dKX�J�j�_���?�{�c^Ս���v�lm7ɲuɷ��� Z1X�?7�]��yh(������[��]�*՗�E�Ue͠Hw*�Z?`����v�=|:%���8%g�w����t������[ݜ��z��
�:�8 R��
C��7�R'��>�zCӼ<ѽ/?O�	|����|��dD6���Ҭ�\N�RW{��-[�Q�e��#����Xё:��M-n��P�!�τ)km�����)��|4V��t