XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���zU�x����E>��<G�ز&t�ܟqј�kXǢɎ�+��Q���B���lZw�����+���	��z~��˷��x��u�Ð��������NG!@ �N�6��0�Nq3{�v�	��\�@�"�x�������X��]j`��X�(:��4bR,�H�5���C��]G0:�&����9f�EM?v��Qe�|y�$"�I5�S;ߤ�f�p'i�O�`�S�S��O`.UWל�����a� <X:h��_�k���n����sY����3��#dj��p� +S��r���k�	���EFr�c?� �@�ݔa�g��c�@[����w�y2ؿj���lY�	��e-���g��;O��m���q μ����g���ڣ/0�Z���}=��&��z��|�^�d[�捠'�b����_1~��&�X�1�=�=~��yrq�G�c�!��1ۚ�#���k��-[*N�&T �@�Î=�|q���3�x�}8���ߕ��duBRU�| i��J/�Wjr��e�A�;�@iv,�,��^Af����G�-*�G!Rv�g��҈܌z ������=��,��Z�m�0=��c⍣�^4x��e��)�{{%(����D3a[�r=PYҗ��%�f"��_���VF6��7����a��r9��?؃P !+��$��(�z��f��ڞ����.�Q&S��gX�r��R��
����{������[��^�L�1�����2���XlxVHYEB    13ba     770�EX�h��$J 6�*u���9!jA�`�)ͪ�{HyW�TL�n�S�^ځhw��a�������^�?�I���xs��D��wH�&�P����H����&7��$#� Ɛ�r���קH6m�y���e�}�h�J�Ω+�v�v�e�!
B�R�՘{A;v$�
	q�y<0M�t(IN��0{��Ō6����,|c!VQc�n�9Wy��'3W���+���w.zv��Ap��r<y��� ��� ���Cꏐ$S_��۰9q{'�C��:�#84d٦�_Q�%�4�囸���,QhGo��{ �����)8�<;�
*�|�nw��L�ӳ��):#��7��`��>��Ѭ���k�M2=��O?���Y�(,Oہ�;q� >}W��xȮ���SCmb�ݪ�3�K3�1B��a"�%g?�fdy��hg֑܈�� �z"��8��
G�(����]�E��ΐ ��V|��l�����?� �����Q���ʸ���lMp=��/]��:���|������7����ƺ��5]����[|\iZK��`�A�����c1vY�����N��d�u�I�'�#����N�h`u��ߩP?�UJ�j�G�V�j{����ǖ��L��J�
�2����5�A��#����[ɽ�{u�j�?D�!�����W8���lF����z�v�P��P��gy���0X�G��Kk�~�ʤ�����ZOΑU���`�`oH��ة~�ҿh���0�nP�u ���^��M�,C��ȱ_Tə�U�&!t��v+���U��ey�U!��WϫTl+<�JΌ���|!ް���� �O�@ :�S�y�J�|� A��K�M�K=��j������$����/�_�i���.�������-W��F��E�.*�dǺle)<�l�T�t�}��0;/]��
��{���N�.���0��LV^�_�s"��\����!�hr߀�]2pYw����&].o��N��v���K苃0�e�������Jf��?�>��}���*x��Q���<�mGz� �s>2U�@ד=����K���!NY��c����q��h���o8�f�8��0�Ƕg�a���S-��7�r��>�A��w�kF�\�I�﫤���ڌ�0솦T5�0!BB�ώ��-k���_���h}���l����Ί�8
��4�Cq(� P���	�Wp��U9Tjߋϊ���R�Z���d'�w���ݩh@���7��>������H��~D�V�5o>�仧,,�C�i,�gv�Sݏ1��H�P�r�]��q�v1�w�{4�H'P,��"��`���l-�
6A�f�0�r��	g"	)
��96�۪�P�h�}f�4O�Pih=��x��IC�>l'�`µ]�I&fq��D����:����ϔN�+$���~ؒ�X:Hs���c�,��4کƸ���p,'���=mέ.�8RҤ� ��������a��c��Nu��l��o�l&��V%����r{5��6�e���k��_���I��{�%o��_�9[:��	Fkn��'c8qs�O��e��<C�W9�Q�u�	�fD�]v?��aN�v�����$���ͻ�=]���D�F���"vbƋ-��/{{	v`��SW��0��2�M�(���G]����@�����K*�Á��C7��;�.����D(�%{fp�1-5�U�^]E�6h�"�$in���줻��94��piQ�Q��r�;�ll�ڋ8�QJ��C��k��GB6��'��4-l@��<`�?<jC�5��gD��.�u��f��u�����_s��	�)�zU闰���\GQ�w^�g^1�}�3X��g�mB�s&��S#,