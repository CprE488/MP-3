XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��PZ�YHK=�$�`환�H,�1Y�⃃��Y�9���o�
�Brf� �q��Y�|�"[�k{��1L$<C������q�����5m/��o�\�N�pRٷ�u���r7��#��)���b��CMs���H|�bK��lR��"C7��Hz۫ƒZ��-�$j��[N ����M�� ���!l���]�s��UñT	~O�q\�-n��^>���}�̀�7�*���V�����%d>�~��ڬ
�0*@5��p~T��l�􀰵#�[tu�٨�X���28���A�{����RCe�T�HXU �	ꚹ�;K�0T�*�����R���TFue��v�������e��5�y�L 3w����j��H:������5@��!ܕZ�m��kÒ��]q�k%Z?�J��^ZQ��Ћ
95L�+�Xłb*@�p�̾e��dvL誣}�0��7����]D�ࠢ΀p�M���n�M�.�x,� �8	�G%v����4���.�Pi�ORFw�t�Q˗�b�I5���}�Ij�D)d�GQ��@i����=��e�#�'T�֛E.e����NKe�,�/�!p��ȠW�y#..GA�Գ}h�G��I��r��H�O���7u�i_k���2�F����!�
6���O�x)lD<}ȼ�2oRI����MA`�E:w�m��vyˬ�H�z�� ^L���EA��~/���������D^���/�|�&�y\1Ct.J"��Nb���G�{�ʺԢ���XlxVHYEB    fa00    2040��K�IJ����V�F���Cʀ��h�!V���qx��1\�Pf�#�LA7C?�ߖ�G�Z���Xǖ�]ݘ�#P�1'&��A~I��)
c�m}#b��G:D�Se�2+���8���w��`��,���*�c�M�8�8�+�����~�迁*:|ڬ3v�n� &Aén
q��EH=�葫�\r�\.�D�*��?4�r��P2k��W[�����R��z��8�J3=g�3򏏅�=\�m���Zz����"K[A�,����a�����Q�Y�]sI�µ�2|.�KII'�y۝8:�5wX�P���SOlD���]�g��j4x$�	C���a<3'���רP��y7W,۞�g�C���>�v������"��1������=)/�}��g�� b��R�	ȉ�_��%��ѷ=�ڂ)
�gF�-E�؇V��� w�'��^�I�/- D�s�F$��{�Ր`��L�E相�m���tٓ�� �5)����-n�;q��C)��7�4g��<�ݓ���k�A�$�Z��\#U��qgʺ/��>w��؆u�������{�����~I���]~i$L=7��h|F�ǡu�{���AZ
���0��[6;�	�*_�#rD}e����h	����^�t��.�b�bjq��8Sr��z�Մ�q�E�X��h�J����]z���!~DF���%L��~�xࠎ�%�&�������U�����($	G�P�Y.-�^�C����uѱ�VC f����SF��Y?�#�-�`�-�u�B�Ú~A���+[NmsU�|�yJ�Y�(�
���A�)�������`fgƒ�oHa���c���g��+���t慍,j��4m)5����~�1f����l3�>�����	��u��6~_�/i.
_���	r*�nֿ��
������@��"$�[F���%�a C[�!�i���}M)�=��.�x������՜C���6��(` �t*��(Ks�77J�#8"���+[/yB:b�b��� As�6�sz8��P1)��x���N��~��t��Y����с���b�tv�jw����&@ Z���kM���;���gVݍ;G#���5m#�3�e?w�sߺ���п�bTI���V�[��0:0���W	 Mm�N�\�9��##�H�= \ҡjDrL���3�>,���;�glLO��@B~�����*�x@����#%��3"�nD"��o�*8�����i\�^6�����8P"���KQ'Խ��[<^�O���ܲ�\��*�/>��/h�*��/o$�6�������8�Vsd�B��y�a�S !�G):�ӽ@�*���"؟ۂ[K�b���G�}��T��i�UL�8����^t`��~�fF%���~�g�*����>�
*�Eٕ:'��W,�2�Y�M���I���g�{P�-G�3(��t�>~��v8D��ƞ����" �DZ 3 Ҧ���˛��J�>Y,9%�qC���0ܖ���j�l]��x�k5�!�B��˴�:@簮��N�|pW���f�����������3	-���dS-��x*�p)��b9R�u��}�������݅�t����f������B)��zm�G�{�h"y{|郸#��)rp(��� ���c�@�Djyᩬ=D��}�ˑ�΅�R ���e��j�j>����߫��-��e=I�К�QI+���.�W?@�:�p�nC3p����*V�$����'$���"�T��堃��ҋO_�N�5Q�1���N��˜���n�����aZ��q���1-3��t`�)(艘q�®{���F1ׄWI,&'���>u]�2���F�~z����:;FyK�<�a2Bz��EѢ�,�ͥ�0k�%z�w�os��1��UEj2�_����N�\�`�CsJў��>��Z��(�L�oB�L�}5�V�X�E�{�8wn��h���%A���/��F��"�(��b�}?�E�-?&K��I8�Y��U)�9*�憵�*u	I�ZH��_a�U��}A�_p�h9����&�?�#R�6��1��G�Ś�d��ШE��p\U��H�8���G`n���^y:�]s�Ԧn�CP��ɭ'�zr�-э�bn�����7��缍�):D�)&H�"\�µ��v���M�GL~������ݮ9�
���p��#f��_PF�A�+��n�?<��rUNj59�J�����5-�w�o%;ג�~��l��0X�C��o��s�j��F�6Nw���G[���/(Nf)���������G/�	PC�v�8�G�L�������(�-Yx2��-3�i)Ҷ�`�{;��`M�j;���I��ﷴF������g��2v��� {]��*U��NR��q�p�|?��hh�~��eC�Q+\���"#>�*��g:~��%��(���X��h���  b�'S�#|_�!{�$������I=e��Ͼ�X�_<F�i�T
�M���!&�jB z~X�c,��>O���9��S]���u`8�hw�k3�*�P���F�i;�Zf�ĵ�b���p?�/�����/
DY��'\��6�s#yZ-���C�k���:e�^�n"_@5��U:f��sΓez�`�mV��R+�9���?>�(��hH$^@�: ��9�R�C�3y'*����Ȯ��ܔ�'m�`ok��d��`2�(��T�ǻPd�f:}��N��x?χ/T�'ԗ�a��5Ȳ�Ycr���:��3ׯ\�-
���A�Ν�1�����5x�3B�9���IZ%+�kF���ph\vem��NF,��C�"�3)�w�:^��@�Ɨ�9�9�x�%��A�Z-�XU��ϻT�~��뮛� N�X��GI�}�UCE*�N�nN��U����NB��iH|�����CM�+P��	Bz�{9�݌����>�4�Yw���GA+��?'K�=�9�0'�L;D0&V��>�k�@25 Ig���
��E�_ab��dG�k�汤�4�i	36��2��qWM�8jZ�#ue����.$+�w�}�%��x+M����I�ᛖ�Yz��q��.lOU*��X���Sn"#���W������VZ]�܉�"[BMU��X5���1��r	��o�0vS�טA�W+t�E��ݯ�W
ַ��@���q���[�P�$2m4�t0���%��+�"&��?�Z��s�X�%�*VB��������5����yX�JK��g�n�q4 ��`ch2xU,G�����SML+7�a��4`?��"��A���[��7��O�Y�!dK�x�Z2�t�9�� (a$��H�e���=#�n$Q�yh
�!ӝ�T¼˜6l7;A��-C�6CC��{E�q���&*�.=�g�_�+%ؚ}�Xe���n�v�S *e���T��eN���9s<���q%��������zah��0�y��RW]����F��77BXTj�wV�`�δ<��BY!��=�����:�)b4�������}x�IaLNL�r�j���L~pB�}ֳ�i�oU����1N�OZ���RZ'��*,�wD���x��XY�,S V�H��������=s�r�4X.�/Ch{.F�B#���򥾃1�x�R�<��;j=)�c�Nː��(%1��8��PWZ�Pj�^�ke��Й.��v�v��&Cb��k�l����E�-#�4�:�0'��`����G�٨�%����v�t�^"s��(=��
�x��9�9v^���{o.����OJ�q74@Ѹ=��	*��稽&���l���������1�_�&�
Q��-?�����4�"� �jy@�Q�N	�;d��M��!�(?�,��H:d1<A�����pA��%b?�XP������l��'？�(:�Hf*c�m6�Sje�0�G �~u'E,6�@�8��W�&RZ��m�Y`w��/MU���* ��U�8��.A��e�Ĳb'�Z���o�͙�7K����]pV$` �Ǡ�!k��D�V��pEP%�q��d3a	F� �F�e�po��H2x�܎3V��.���Fu�kx�չ/F����%�\�M�j�g�c�U��UbL�q�l~7��6h�eۚ��x���U8��y�l�s���ơ�Y�N�Ͱi��D�h[�8�68��p{����*����q1�i����@�~',n�8�\�$c�_�ul����o?��� $m|2�'a~�yyi+��#���N��l�pj�(�!N_�$�2��9�M�%�7]tL���wvL.�����Jo�A�����'�u���\Q�T��5��KNp
;���q{��˘���ֆ�f�k���1g����=[�{1~��o��cf!ɨ�TIļ ����E���3�7��y��eڭ�D2~�x�u���ʋ�,P��e�Ԣ���F�m�(�ҁ����hiEސ^����ʶ�E���#��I��`닜�㹆TOb1�l������7�XRχӤ� ���<�Yƭ�$�!���|Gp��:'Sl�*���<s&(r�� �8�Qh"R���d8*.q��N���`��
�d��0,j*.����Z���7cϝ<G�r��tV�;8�1��|T�M�"����AgoMQm��&B��B�F�LA�ST6�cz��5���CЩj$��1o��ή��2R�a�0���>�ә�B�F?u��ˆ���WUe��"w�{����X����yVD�$a`����NǍ�����6㘀Ig6={\,;�Z��/�v����v�܉좯*���������lZ���\���Ѻ�ԃz�]fȹ�|�|^�=q+|R�1�فW�*agѧ�9�f�n�x�3�?Ϯ���/��k������H����g�d�y�|r�5���r��/2�9^j�����]Pi~�g��?��%�`S0��1Ȓ�\�b;�����;�`ط�����0U���E���Srcì
��#��%�Z�_���#���!���)p�S��d4�,��4��l����䱌H�"nƄ	�|�5�7TM���U�#�2�������O���}���T�35>�*��������!�t���������5+1���hJ'�����K�ꫯ}h�����U�#�T���(�r7�{#M��g�J��7�QNm�7n����ꃛU���G�|s�2w���$����\�%x���jo�ĮK��^��k����kP1$ �w:Q�v���W`�l�xa�kA�����N{<����1`�u�o�
����#��7C��C'`�C�b��	4��f�F����C��2�L��(j��x6SAN�'��"��۹�H�C�ݖ<Xϟ5�I�c��B>��cP�9D
��k�0¸џ�ý"5�.���NO������A9�ž*A�$���
�Fa2P�e�/�������V�y���&P����S��l~E��ت���*2��NoZT�|S����}w%8���f��Z�:rZ�n���}�&f�ך"i�nd���
�zqڢ�C�&Q+�WF����������0>�?��;�fռq�s�����c�_�j��l�&));:VpEN��%�J�sa����W[���*%j�)��A��H�h��o�^�(8��[ge���6I>aR��`X;�\���ߍZ]ʫ<o���)׍�X�@ ��K���,���NbՄ���!��iԈ�Kl�.�$�cC�"4�\�U�W���i;=R���d+���`m3G�5�ܛ���2�ߟ�+�	�5YO�{J�R�����K0:'���T�K����o���gE�Q��X���r�Dغ��0Ұ�P���W��o�9�� �љjՄ�M�CȘ�hL��HR��vV�{����?op����Hׁ��`H�l$����;�U|��Cƃ�݈����v`�Z�^��M1��
�mP�hê���[�x$.nEL��ʮ���+���LRWJh�z��������D��Q=��-_�����<�y�R�hʹ��so���YzD=�U ������*�6+�\�^�vy���z�i1��+�$_'.��X��m*�$dtZ�i�*�9K9#�R��9�Q��59rt����ڃ��gB���%d�N#ݧ�W����t%�&D�r���i��ȗt7g�;@�	M�F1vw���P��2o*�Kvd�.��khv��"+rT��mR�������P�6|;��}1Fg�;�l��W����L�����Q��o'b�%?Axq;D߭"����mA�j�}�(L��������Y:8�U=��U�	3�w�����[E�&�pܒb%�(ϾO��^�2��^@�rد� 6;v1%���Uu�ؐqUm�W�Br90�Mt;���#a��ف����=Aã[��2��liÍ����Uw��¤��e��_n�@J�1�_�_���j�f=�ǭmJK��<D��}�YG6F��q6g�}��
7�Χ<r ��rT�\\z{x�����!Iv�}p��(�L��KC�Ho�a���;�)8��}���z�!3P��~�i�����r�A�<������MC'Ԑ�Z��8
��$�|ˈ����y�{�K�W�˯�
�OF�M��>1���ȃ�$���ɭ�⊈�sh���+�Vut�|"���)��k�c]�}�b牉Y�\m�th8��v�Vত���BB!E:��~B[���yR6LAc�Xz�|B(����Ǆc����_`�_ˤV�p4��o��������v3��Q�K��l~W��vF�)Cm�Z�Ffk�?O"{�P���LUI�W�<<����
�7y滒�}H�
�p��5��"��Ҷ�gdG��n/ �5 �N���u���m܅��©�O�i��m,�j�9�y"�Z�$jLG��q�yā2;ZkaW�X�7�D�8����1'Wû'�m�i[^8sl�=��:�����|��s�"0��핒V��;H@�QE/��Y��^�gT!ZG�pA`�v��n�P^�\�����纺#mDM�����P��<���X���D8���-2Z�[��t&|9��֪�O�	.
�1�ۓ)ƒ��I�@�}o�[5o?(q� �C�X�V3�~�V-���ᩯ,�G4H�?����D�	4gD�z����\��{�V��:ey4]mA`?�t�0-��˘�x�� d1)� �h�+lv���ә�$���aח�ވ�a;o�L唗Q�z�ct�)��g��J`�b��n)b����-����ɨvW&1��I�u�p0c��+΄�R,fɠˋ�
��q*���.R���n	�Dڮ`1�z�W��[� 0e~Eo�Z:/�r�ψ����X��������4��A�u������R"��KL��,c�(.�w�x��X�}�o@I�1h�e��{
X�p�8"#k�#8.C�t^�pgC�h�(��$���LԥȊ����b8�oCJ8����+�\iB�����"��AZ$���V�]j� ]��a���sl?��ϴ^
6R(>�@�Y�^��?3��λ⿛�>�	+�	 e�Pތ/���;W"�`�V�W�(q��0ܟʶ�����0T��*�\���pى鼉�v���>�z*KQG30����K�.a�ԧ��Ʌ�Q�+2-] �Z�hT�Y)V�B-�R��ʅ�{��U¬����$�d���ɘg`}1�XQ\�a�m������?��#�c�(�i�)L�3���jO�:H�÷5���C�J����48QT���'��	����M����شk��f��s�W��H֞j�l�fu����n��3�m�/lu8��i���?�f���,��F�%O���P4ʼ,����	�!tNG�����)�Zz���k�{^�M�r�Bf���%MB���XZ�,fl�����%e�>)�/W��a3��0ntT��~���\?��i���c�`�%'�����J��3u����g�{9Jn>�؋�&�AEyv�j�;�z)^����4~B
 x���2�lx����
���(���W`3��:��G.%�L ��'�]�g��&9���T�����4��#3���g�j3 g�7i�z��KH����C���҃꼕ϱz�sx2�{��B)��Ɲp�Aq�֚2O��)K�l�� ��&j�x��1xmܢXlxVHYEB    4f62     b50�ñ�З���iD*��>TO�ɲ�%dV��[�YX`��e-�B۾��fWӗd�mHܹC�JJ/�W xDm�J��D�r�$��^��K)�i��&C�b�B%7�X�&�(�Qo����!gr�:=o��*@�̏�pB �7v�̽��R�������
.�i�X���ᙯ�!��+����Eĭ�GfYgC��%��m�Z�o�sYY� TT��j�<��A	ϏK .Ҩ�t��φyhUN)�|g0ٗ!~�H�5��)�� 9^�7a��yh�Q_d�Yq��ʥ�0Ji��� Յ���;�49ࡓU����;KQ���"�(����~��É�"W���~_���'g}�;r����%S��	$�;��	�y�'X5g=̄ȣu5v߬�+�FZ�� �9�.�Z&�b��7Q^H("0f�����S,]��o¬_?��o��A�b)�d���F�M�~�2���<Sq	kM��%l�ཛ;�vфl�����3sz����걣\r���u�WA*X�$l�ʫ��$êt��MF��o�@ w��&�:RH�s���Nq�'=��K�_�U.��S.RW>B�.��5JW�5�dB��?�Xx%�je6OD��Y�'��� $Ċ�j���MZ�Е��HҚ�!q��[P��5�H5h#���d�d-Q�6�_���+}����RC. a�x�����$��ܯ'䣸�#h۸j��9,J��sc~uf6�A���b|�e����Ca҂�9c��`)�E&?�&_d�;	o�U����'�����q�#��/�p����%��|�WmE�G��<��#���Tyf��1S�Ƹ`A�}���u%�:?�)���2����]`��G�^h����:�6��1�n����,1������= H�}���*��\�Jh&�[�����"�S�㊜�p�>�'gl�A�p�Fyp�s7^��ǮxJ�o`揥�|l'������Y��Pݬ!.�G�!e�KqD�� ��[\����T�ӟ+_XsC)�<l$6upF�N�؋O���p?`�3�~�m
����|D����6��ǲj��#�?,.
d�Ve�ĉ�pV�b���)M��h��	f�;�8�. ��n���@�)h����`&�Z�7d�F3���|Mkّ/�CMmh6�D���V$~�0�����A6�¨S#�M_�I����39���)Ϊ=��d�Z.�'P"�I#�-�L��I��|ֶog�'�nw����\�
���w�7��]}�<�����	T��[A�C���S�h9���lk�╯���J���Fٱ&�)���~?k]�|-��_�˩b�����N�����ȗ5U�'Se��D$y4�MdJP̭$RwڗgO����Y�∼�|�|ؘ���\d<����L�n���O�ڎ�R��k%�z���-��������@i9b�6ɗ3����O=#>-�W^�i���)�����3+Hd&�sv�T�����HB)�4 oQ+�M!�b��{~F� k���\X�"�/8�%��%����	8��
����K
-�/*�v��q�Y~�Sʆ�H)t��;L���������Ow�I2A)q?M.*��@�|�2���Z_��d���˹Pmo�j����)W�s�q�����q�𩕦F��X�Ⰿ�WUZ�4�EEK6����g`F���H�������2	��)KhM�D�-����E���#�4���)ԾŲ��I�ؐ5�'��=_<�G��J�R�H�臀@�S�7�o�[�m��R�rO[x�@ZV5ͽf�hQZ��D�=&y���"�'<��"C
�`?��I2��Jtsv֓����g��pd���w=z�r�'�$on�p��M=��kO�@�o�a���ƨ�ES�;�'�h�]�Ɵ}��t������uxmlB"c�ʴ��J/�{v�i<����J&�%D�g��t:���Pk��B��D�&��
��w�=]K���]�7L�<�i�-�?l��7 �OB}�h���Ʈ'�e3���k���~b�v�lx �x�E�E�81$7,�Y(��'��
ey�}K=���Zlf���?�{lƍ��$��BX��1Cl$-�Ռ���Gگ��R������1(}�1��#ď7ցL��Q��/ǥ��Bv'3�B���,�ϲ��MjwؽEg���A"����t��M�H�޶�d6�l���i�ZD��$�������B"hm/����Ә9�3�����$ba��6��1^�y~|��{�V�*�e��� y�g�[j4܈��k�5u3Q��J�F�SbQS�/�u�R���� �3.�j��E�/�ي�xcU�k�VDv��J��4yڕl2˴I?0A���6����Jf	�"~����:����t�#�i�	��<@���Y;C���}�y4�}�����vS��)�GA��x�H��!�1{n=u�Y�%Y数��Jp��np�ވң�Cz�����#F5���'�!��/�6	�%r���3�,$Sٙ{�yu'��;���+|�֓�Yu����jnN4��9�i.�7��*��dKp�r���B��~*���1	��I��Ѹ�1��<��G�{�A0�h���ao�(�X�`�Cz�&���{�V"�--�;$C]8��׷��_L�(ij `��3��c/m��&�%�mM�I�0%,e�7�.B��n�:(�p�Kz�������E���Tvb+f�)�9�'<7�^��'����onk�l%��jq��,۠����?yam!q��'��L��![m��Щ�U�9�2�����V��7=����cz���h��k������V�K�G��+Jc���co'N���NDla�