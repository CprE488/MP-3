XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��AT	�)@����!�-��^�8*"n�,Q[U�Kr��#K�}��Lj�����_�R�m�?B�%�2~���.@[X4O�R��TW
E4$�[R��I��e4o���%�9=��Ƌ��%Kh]�$g���^ϘN�H�x݆��<���F��\���}������m���n$c̹t+���oL^Mܘx!=�n�3�B�e�c��њ|5��U��^2m-Lq��Om�F�P���d3'����!�<TT�����ѓ�P�/K0�!cx5)(��Рy�wW�.�\���(e4����_���G�>m�ŉ5�z}_~�.d��9�Sa���7/��ћJ3Ú�&|&'CSD��*�������%l���x-{��5d`�K�E�����o{9<��w�D��Ҷ3���k���������P�%�f�>�r�$�j��r*�`��/\��&��*�����^1�_t�Zv&�:�+X���<�ts��<��c�)Hf|S<�n9~�1��r��h�g��Me1�I����
/��zI���H%���B��kS������Y\k�������&��-5&u֞�[����Q�l�#[k�g��DS���5�Vm��2]�.�a9gh��R�5�iq��&a�$�F�K²���6~��9��?A��5ˤ��[:n�b���V�6&H�X�x��N���t��՘�Pxԥ+6�ЩN� n"��X:k�c����6o;��6���r��J&��+�K�3Y;�{����q^����XlxVHYEB    2b39     b10��q�鵨�1(�a_\o�:��_�;4.T)�b��^�+�}OgL7��i����������8�o�6#+ڟX�Kg��#�I�A��HB(4�����ߨ�Z���+�%�������� ���q���_���ZE�M�#h�KC�V<_��bY�Zp�yLca9#P>y�*�}�j��:��c�K�~[b:�L鍎�H�m�Գ�O�bMOY�qn|��@ SSL���)���YhB�$���p\��N�}�r����_���B����;ϸ�%L�m�\r�^S�� q�"�3� ����1Z�u���H���V_Ot#�ȳ�r��\ �a?���^ODe������cB
���v,�x�v��T4�$xD�!���3�|Pլ�ӯ3�C��^B��"�W�gzQ�<J����*���'m���yP�����k��^-o��*U}g��$�fia��nw|��#fO������I0������'�ܜʣ��97ʸ*#�]_uT�gg`�����¬� ��I	 ���7U<�t6k��>O�������tHyk[�T'(�+]���r#�pk�g�v5�#��Z��}�mj���â��9'�o�0#cFC��i0j2U�[�86mQ$]l���ȢI�W5��xS��|/S%
`�<
4;}���4$#���V(�t@�At��e��M��s�F�z�*@�^��M���V��i��l�r�6�y�RA*�lF�9/�X��O�3��LY:�+r�/V��r���Aj�N[ܜ[U����
��9�?�\�,��n��Ul��Uk�ڝ[�oE�mǱ=�[q�A͕~,�	����/��=��!�'�M,'��ؖV��N^�nm������2�����ם��E�r�(�����i�Am���N�XT��Ʒ���xi`W��e`ϴR�./�)���w¹��/B)��[��=T$~B4�T��{@�ozc��#A��5Qd��L��8�?�ahQ[�m&6��S|Z,�Ż���X���g�fQ�R2����Q�p�샙�#����6�&��s��Y?��1�_�¶�m�7I��H�ܲ����)&Zhi��䴙�%�*��9Io����pt/_��a�����%:��AHik�Z��P:xM�%}�CZ��y���Ӎ{�yA�郞�	�Y����.!�38��ɀ�|�Ɋ����ھs̭gfQ9��8��Z�uU��(�-n���޼�&y9.����B�s�kD�;�D}V�o�{��mW1�Dy�j�ɟ@��Ze;c��fl���r� �$!�gҌ2�����5K�_���e3m��Ω/�P�l�]&�������*r�e�`,>��:f8H�L�Ow�x����~UG _��}:����z;�Tg%�\�KVVLN��K)��������k'W��0z�![C՜�dpXf�<('!"���� �!���\2�Q�=�1��̗�0-�]̇/M�,�i*�B�����t;a��r��;v�/?�qA�2`M8�h���I0��w$���u��%��I��ȩ�ы�*�ڵb�(�V;2���I{L�k�֙�r|J/�K?Dz��d��l�ώI�8IM�50#�-��M̄6�&�o5AB�o���k=��,E�Ϣp}J2�B��wh��I��3���
�G�IO�g7�UhB~'z�d��TW��8��)��f�����}�~���\h�IpPP��a�nU����M�$�J4���Ī,J����яN�A��:7ň+-�$�A��~����(�m�:�(v6[Ԩ�C^H-S��;;�Q����BTqx����a����q�̖m���g���[�e���dg~kƧq�	"
�x~���,;��li��<������/m�a�	�Z1�W^����Q];>�
�|�����C��̲�9��؃�,��'��o[�Żތ�E�1r�n��M�e1�މ!��]|"��(�	��tጃs��P�����^�c��`�،������&c�i!I�@UCj�{�K3�ص�����F����p�\�!J�{�$�\��:"�>�(ؠf��f���Ɖ�
�������G)=���C���'�#�F5�6��ڴa�=k����]DJvC��L�w�����T�&
z�_��HY�lUx$�J�i �|�;�����{��}�_6lr���7En���j}�,62���I0�I��%Տ �W��'�)^�W;V	�gW����
�B�� \���<�ny��Eld{Q��t�(k��"��B6#��E,�g��b0����rKKY+z��[������#i͠H��P�p��!�HXRc`R�>�����ת�һ>)O�i�sy?�� E
$�]��˧���H�!w�4zNJ� �bC;04�Nfz�%����C)���eE �L[��΍�.�=W%�����]n�I��ޖ����;�ɩ5����I ���H�F&�T�i��m�"5HV���5秮�0��e��K�9L��H�jؓ#�I���~24�� z$;s�O�స�c����"�����HJZ=\�	y��SA�U��"�=l&\9/M�����2�8@�FN���Cz70fN.f�J�UV�ĕ�>��k:���.�=��x3ǃ���|�+Ṛ��Sݔ�3{�ܕ��i3�mx�^��D�����L+c�ܒ���ܝ���:�*�Ǚp�<�|,V~('81a��gz�=��)�S1�4��R�~^��7���K.K�%�kb�h�����S�I�>��Ӻ��]���%�����d�o,������l�������S�t