XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��oM��[��5���'H@�s֠���k���qz�Oi�j7���TV��+A��6�`l0EK�\cQu�7����Cw�����ԽW̋�Y�WA����#OR���b��5C�\
������\��j���g���9���j�I����7�Ҧ9��8�D:���U��T���h��=e����ًHM��3k��u�|���.f*���B��=c�[�ܔ��X��&�n?D+Ui���V�����%��<���ki�+a׷v.r;/��!H5ž
�j��F��<�?Y�Pꂚ��s?�)�H�q�S�N�Z��?�*O=��7_Z�T�#Xᝠ��=��	�T��_��흮;��H���Ǟ�h���^by��	��%� ^��J�L�%��B�k9�K5�����<Gw��Z�2��A(bk���0�Q]�v
����͟��ɬ�	C��1��$�Ez�R8GiS�f������W������+��=���c���.
�Ц	:�_� ����k�%CҪ���]nk��������@~��;���l���#�t���D�Zpu&;��ЙDw*D��}��͒j��x1�w�
>��j #<L�In2�W����}��P#��w�n�����@`
j|��'�l}�1���q:��ڥ&�_��=$�*�_�+ܻ�r����c�M0�5�h�He������U�r�����?�[i3�P$�n�T�y��̤�!�5
/��70��OT@Ae:�a.`?XlxVHYEB    5866    1100ǋ����:���o�)��q[0i�ױ�L;M����䐺��>H�X����:�nq��+ܳv�>m�����Oً���'N���&��S6
�<~Wy��4J�x\��\�&D5��J�?EJ����6�����2Ym	iRM\�f|�����?s�??�)2��7h�����c�-C���\JD���?��_A�d�T*�#`�Vԇ�)£��D�K���q��6Y�j1��/��O>N�p~�a�H�� o�B0&��5!v&�8��l��C�/F�?L/ڑ��*׳ f"�ȕc�1����>�ھօ�$9"��9+ 2@�6�'��Y��$wOp(e���X0h�/��/�]}E�,!��9���T^��HE����4Cj�/��z��}�S�UayC��Z�vĥ�����'��^f�V�_����gA���ɺ��/��r�����%E�|���큉Le����� �U��\M̼�%0	 u&YΒ(�"Hl\�&��h��J~=��z��<Q�j���e�j��2:�ґI�~��7���=9��{]�|m�~ ��O�'~���"uu=$��Gk)�NZ�D�|�b/�s�Mv+�� �2��ŷ��V&ݬ���!
����n	k�\+W�0��������d���'e>űc��<�`���=����Ծ�W@���>�7�f�����d���a��c�x��bF��_<d����{�]�����*0RL����2�̢c�zj#;�5s�&�sQR��K���=�>�9F-��Z�׌T�]��>hvO���B� q��}�pHTh�nmSu:Ò7}�^E�Q3O��_��ѹy�#<�*[��
Z*5V�(��!��)�{�Ox���2v���M@��_f��&��~�A֓(�e�ЀrMn"�M�ݯ[S��&$�������kv8�������0�fp�o�q�-=�'��`���5r��V'�I�f�S=y+�26ͭ#������I�%�e�����;�����{ݧ�@��H�p1Ρ�3;���ۄ�7(���ԥ��E$9��:��u��R�j! �BDhT�l�$G���^gr�h�;���O��}a��v�������G������t���ׇ�E�Pk%{y=#�D��Q�'�v"�#z�Z~�2!���%�z��i��Y����9֞t����+bK%�_s�Ĩ9�o9�� M+W�vaX�0��^�I]$8�D��M<����q�?��4Ft�=��Y̒�ӯ���y�᳑�jzJ��!%8sN� ��t|�|"�A�����]�p�^C�M	����1'C�`pY���}S���Ĥh��@���	�Z�в_i�	��d�vTp�v|�c
$֦O�*��#_��K�:�vx��O��*�����Cb_��,g�xf)6�0�4�?4����= Y#,e���ik���slGε0G��f���CE���hS��@�r������P�\��V�ĭ�B��v����������!�Q?�Ͷ��Ѻ�$!0pN��(vn8�����%O	� ���8��_�3l�o�a pAUT���}�T�z�a�wly� 4c8-T�%�K�V�/S��q�����oC4�S?fFi@��r��I��.��Y���E � �i���8�����!�
h���B��.�Ub���Ԥ�S9`Oh]�?]ĝ������ T�`��;�9
��Α���~ؖ��O���x	 �O���@��ӊ4�� ��6n�OA�����q���������i4��B��d��Ws����,�Bl��'iT���4�x,��ދ�{ў�֌�&��2��'���w��7�̩O�^�#�	I�2�	Q������m��5�E^"��b�/�c8tD���&�u�t ��nC?�YU֌��i��.w��q�i34'ӊ3��~�VS�-��2Tm�ʬU#�bK��T��b@7�X��N��dopSa��`�"����X�۲&n�~�;�js�Qw9?�yA>�H��!�s�q�4�Ƌ��l�hD�;77�#�P].��fH�n��{��	T���/�mS���*���i�2��/��Ϝ�Y��J�X�_��F:��ҹ�٥PPލ�*�"�����;;eov;@���4Ro���w0�)2}����9��`�T�XgH� PMd5�(�C�������D��w/��Ʉr1_��a�JVF��V1\&ye��8�Cc�MJ��>����<?b�I�j_4�x+���D�J�;�`/���f��>��l�a���_�(,�Sb:�d����#���\�8���(�̵�� \��n����j-|�K��F�W��o���q'�y�,&x ȝc��S�(vٴn��óDC�GV�;�����F�SF��"�>I�M˼���v9�)�R�9<\�&���co��z����{_8^��z�>rb�d6j�rc,ή�Ԗ�#�oC@���`��6�
2:��=��Hr�k{�=;��9Q�bH�X�"6�?oX#Y��5��Ęа���h���E�� ���f�+P�<�,L@.��~�9߫���)��)����}�z�}ig���צMq�"�K�(�<��E�����=���|�F�\v�-�ˢf����l异���7�����tC"�߹2:��H����s�7A���G�w��������ӑ������S?��:)A��#�*�9Ɨ�/�,~�!C%���G;�1^�������8�] ~�
,@b�l�NU�Sp�7����FL�_+Y���W�Ԥ�d�NZ�WÃ�/�y�e��cS.�"5j�h\�.i)�fO'pG�J)/�K�|݆]ОM��	��zK<�z�S�M�Pb�!n$��[�P̬������Џ	� O� �$�.�v2dZFſ8� C�`��љ��(�|��.9���k��u>�n_e�������M%_\T�u�uG��j�CД�2k�����Cԣ��}�����=��G�+���D�]F<,���vU� s*ћBFp56ܣ��1$���p�C��]]��u]�����>��T}��H��t�E��B��E�dsaTwr"+^l޻�ڮ�����5[�%}�Ĺz��"C�ф�s4D�ڢ�/�(��&b�g�K�'�������/r����w�2L��\�����P�����:�̤�t8���-�0�G�7��_����rݠ�,B�q���u<ѵ�&�%/���1]|q���Y�&�g��)�ӕ�d���^�XS}�\��Qz��l�qk��i$%�ʈ������C��]�HT�D)'���m����,�ZI+�+�2�t��-�έ���e�jWƷy��A^>����%=J�I#�R�������x�OΗE`as�����0b���&��k	�f�,�ҹ��ۺ�Ec���nj%�@C���iW\���F8�I�ԤLa���bw��$��k�D=�+���2|�S�&�D� ����q��d:�8���u�J5�b&Q����<l�.x�����s��ԋ�o ��%U��_�%����PĐH}Q9%7�N�1�M���(�� �k@iN�$k��p�bT�;	�Ox�Ng����8[gO�H"3O	mKY�)���ܒ����i��ޠ7�!ܹ��{�sf���g�'����������I����$�m�\i�*��z7�e�DjY��*�$����۽�*!YAٗ!�ǌ��5�;�LT��Z��f����Q����hl�G�=��Q�?�c�'�� ��	�|if꘵�Ij�-d�a�R�94���k�A�F'��N�>�8��*���#2�>*k{VLïr>3��x-r	�����A{�>�nK�Y�MG���,����+)�Y����O@a�	����HVl�q�t���(�=����G� :MXɊ��H*[L���)��Dz��6��Ԗ�����N����)r����YE�t|	(��3���(�Yycm�92&#M�&�Jq�<^Г���{��!D�^���j�j������c�bEJ �G��6N�Ù��O/+���T���d?k��2��?'�#Õ�ض�v�i�[�8v�n�,A/3?�$E&���otb���3�w%պ�H8�Ν�JܒSms�)Ī61 5��U	��?ā���~��]�,�6G��OR�I�{�}�Ɂ+Q�(ӻ!���/-�ڎ�[6E"J��-�����N�s��<���JA�����$��՞�������{����l��hؑsgR�E����T��`���>��w.61'��k