XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���w�)h�٥v?�;Sxd�fk�Qk]��R�!��rB��*���&}�Q�����S}'0%��j�?��#Fq��ꋓ^6qxH�L����r�l2�(	���L/?����A��J���p6w�bG�
���ޢ|q����3k��X����4}j�.�4����9A���\+Za0[��VT��xJ�o����iQ)u�:˝�d��hZ�<KɁ0HǠؿI�Pj� ������J���;���H�+��Gv�gF �#���#�k�,�Ps�@��}��'�P��`Ё�b��@|�!L9H;S��4�}-I�Ic�4�>�7RS����,yy��to��!A`�=��e�% |V�� -xtڳ�z�N=M~������HꦀW�-����!�\�h�AWg�u��g����J#NE��8NA��v�[�Ǒ�+�������Q���ο0b+�#�O��6�m@�}ɻ@[#�T�?�����{�gpu�I�M<���mV=Id
D����:#d�3�������
k?B{�6�1Sm�ܾ���x��7D� ?jЌ����[��t��?���Y��7�d�X�Z4�k²� 0�C��E�-V�RqH��7x�r�#�]�����N�I8������A��G;�s�k���Q1�*��W����k@!�-�:[{�0a��is^�
�^���}~��W��sBI�N�����+h"���<�v8~|��"�	�F�o�OS4��8����
^�ݧk�XlxVHYEB    af5c    1ad0�?���K�P���dOߝ%�duG���л\�Z⁅���.��h����!0�k[�W����l���
�s�B��},�Ck��;<x��[x���@�/�{�����^{&�:���pI�����:���s;�\b�a�N?��J>���rd���:"*_�� ��6��%�k����Uw�:v�j��ꮇ��u�7�+�@�Gfx$j+GMh�K��IX��KxKH1��V���F�k^W*������V$�c��oz�HpjZ�o�����W�������̰�!�/H����R���-�3k�/=V�X.S��@��;��q���+�,���X��u.sUdlGN�xu{�a���}�"���քW�D�Z~�I�8vP ���ɨ��½{ӂ���`&S�v�_������$�b�T,HӞp/V��h��/�Zo�	b�I���[�;NGx��n��q-7j�z�-;Y��HY�4H���ȢUXP֢��[�~`E�x�]�oi@¹�c"���@�1e����Xv6i�sk���7F�X�W��7�mHŢ��#U� �4l�T�%
	���uD�<pjKO8x݁�������LgWՎ��b 6���R���P����IH�a>����w��=�
f̨�� �Ơ5��.BD#�vLa�V�l��p_E
<��ƘZ�Ho�g_�F�VV�s��3lEӁ@
�<�f)�g8�F�AB����D���2�(���2���S����(��[�`b�����O謴��h��B��A41�%ҒM�����L�ɲ���q9������E5�º�3)�DpXv-Wid1]��:���H�I+<f8�"�p�B������E�����R�"m�9�6������x���o������VZ���
*ۋ�S�{4r��jP��]�b.�bs�a�=��;]=5B�,kI
�
���󶶤i���N�N��u��S���Dذ2���"8X�Ev@6��Cn�b;\<xG�����}˗kJ	8<��ۖ�D��y�Q�8wQkF�Ų���_��c��愷6͓(�:0,�ۑ�*2уa���O� f6�B!����:�#�y�p�;1���  ���*�Jo�B��,�t���7U���ox�� Rl�ݮ��{;C� ��3H@��b�#l�k��O��ˎam�l\���@��0���E8�MY�s����[i�d��~2$����a�zz�FJ�/�xb,��=�Ⱥ������I�X�Ok"��rN]�6�����T�o�]�)���/�q;���P�S3�Z�GK3nvx,��.�.��x2�p��Y�\)|�@��� Xj4��U2C�ܧB�e���w��{bT�e�Xb�3�N�����z[^����U���"��bٻ@Y�?(�4䲟y�
P�����G?H�����1-5�_����&�J��E�!ÝI����
�Y��LL�7�,��ÓT�$���{^������������b&fØ�Þ�-��b]5����c�w[Ӣ�ނRm��~?����UWȱ��H$��h��F�Ti��Ϡ-�y�gď.�Hvi4��j5���T/Z�0o�]�V�N�:�q���n��߸���e܎�������+7|"d��G�&��hk^�N���Yį�j�����}u�םG3���XD\��}��ʞ�G�32~�����vx��ɛ8Ba�"N���2\���0�p�	49���a&N�V�s1�3��>�K{�+JfIpY�T$*�Uԓ�"�J����O�;��Z���,f\	��J��ha웪%܊��UAV[
�JK94��J�ܬKS�#�6��V�5t�� jP����ƚ��� �6�_�>����=�xh�{N֢�&MV^����c� �]�ZKp	%�=�$����Ӈ��+E{�-��jܒz��X��T*BU#�[�I����>��S��i�%F���g�f+yo�g���2�m�}�~]FY��[����O�3�dqd�[(\z��y����N�`| 6@�����_�FO]��J�N�$��8m��`_߁��<~��@
5� �ML�� aw�
���[9.��j������fu�Ba�Xq3ƌ�L�Rي���q�_v�GDW����G-@R+�D�?��]��MV��|\��_�F����܂ֿ-omf��R�E�2)���J�IǑ����B�ǝ���M/
����d)�@��a�!v��Byc��O'мi����q��)A^y۲��)=|�j���Ļ�7=	�	]Z�!�1E"�l��JۅB,��+#&w*0�ђ����S����d�)�)?j� �;�-d�mɉ��\f��@�17/T�+ ���FN�$�D���R�s�� t:�|�!�a���c̽Nb�x�%N��c}ݘ{�9ܒb�����!�䔧KXߌ�m\o'5%?���N����amT�7�.D�ԟ/�ʽ,[y3?g��}�Uڴ0��QTSŮͻ2Y�i���S��.�VXПS�Eq�́��;8��5]%�������;x�)XY9�q�L�1߹��D6���p#8�����,nC�M�{��)D����SBF��k=6�8���'��[Ɲ�5DG*B%��Wai� ���{��7"��Lx�)��j�U�.��?� P9\I>�X���R�b�OO��(���;��?�sG��+A�9��)���6�� F� ��Njm|e�0$胕=pߛ��H�{\���ʳ�C	�܄_A��6��1?�O����"��K猅�P�-Ȝ�п��\)���o� "�5u�m���{$>J�(���`�"��N;`m ��8	!�c�4롑��a���XkLw�!�E=L�l���G
ET��^�,&�E����� �sd婔`���e�ϫ�AP���ޙz�ɸd��g�� 7���I顬wJHڦI��P��?� r���k-���D��jeO"Ǒ�I�z�A�Ѫ���	�3�g_���V�k� _yt@������H����R@$��M;��?| >���Sd�.�~��뇏
܍��(M���i�b��X�ͼ,�;��R�2�w��9Im�()~��4Zp.�s)MT��l3e�*��ߟ���Y�t5�U��q�g���Q��J�[[�HN�_�@H��^Lp� kz�E1]a�A%��|sKL��82���Zl�X�I���1d`���s[)hݥƜ��	P7=�b-5��1��b N�߂�m��O����E-����L�I/�������g6�c�D)O�@����0�-Rd}�����T�H�p�Ok��N�j�G+0�P���x����6�U�r~��!����'h���%e{Ɋ���'��q@n?r�i�L˶��~��G]�>��
�:��>O���S�L�9�X�j~� %	���m����3~�A������������=�ޏ�~of�/lv�c~��	��0��\(Eȱ!�n��-��3@�&��V-�u;Dl���B���tC���؉b.�������� /P�K��U?fݑ�ϗ�q휕��I��{1Y��c�)��C�kdZ��Ul�4٣��]��Ɲ7
��l�x.�B�*S�Z&^B$���#������Lv���2!ő
�_�v��;΂��%�3tu*��������	��-v��S'��H��"z˲{|�ڇ�_��b>����v����>塆�kYZ�z�tY�=+I����~�gbA����̣���kVz�X�Ҡ�IJo��`�:�ȗ�B��\T���ʢ9��1�����9'�G�i��K�+�#z\�&B��L�$B|9Ѫ��)a����6��xc)9s��\�p�:���"�yU�N������np%�I�b�F8G~��(�^�m�c�d�!�����(u��t�\F��qO�y�._;�a��Y�2
��;��EX�>L�1�O�ɾ�<^T�enR��Ns o��'�w{��DJ�`]�&*2)O��x)e�V��#��������pы� hǍ�쾰�E�;�⟗}�S��L7#�Z��H�'e��l���*'��^#P�C�$~k���	I��[�תU���Y��(ꔗ�%	f 9p��<����2����f+.��AD^P_��Ĳ�;��iw|z&�yݶԪw�[�Ux�Ѐ��v�_�Ӛos�c��_�-?<G��tPgPv�UsV��� Z�!�at۾����٤���r�]lܘp���sg���� �(i;4jZ��/����=b��Oa��jXP6��g����b!Z9`\C)�>S.�C��uh�����-�l0~*����b��t}Bդ��2,� �۟��	Rnn uE8X��e�Ƿ}7����}�#�{R̦o���Q�I4YWȏ�� �5������	���M����qC'^�l�h��R<�e��Y%�l5�y<|j�uJƪ�AcI#�J�(�z��p��Ow�Vg �̈%�la��UR�3�T"n�OwA�u(@��M�����-�����ca�?���wMǘ�ob�|{`j�|>E$�j�!� ���\M�&����,�����S�e�3]��1�e:����E�7�ll��+�������`9����'%��qxu��ӘN1�ie��*>�W��1��Բ;2�X�����Y�@�ׄ[�Xi4���V�g��W;$�L/4-13���e�E�0�c���?�>n����v"鄉��U�9բr����5vj:���F�ү��<�_��N�e7BlT��f�?�R$��S�$���6���p���JCG�z�c����!w�Lɼf�­�K�Mh��g���z�n�h[R]��="��%���;ɘ���Ct�*\;ؐ�S0��/�S$���i6�F��0jÙ�|�~L��2R��L��
TVA�Z�*jh�b4M�,�~�4�l�S�,����b 0\�9_)��=9 ���m��lg�_9�Ì�i'�6����d'�m$�X��4��#<+���K�D�z�Θ��]xI�yփ���>HJ��>U���/����/�&Uf�v9i�i���M��q}�N�\(��!_�\�Mܱ<�>��'!�N�u��_Wj�?KK5�##x#&�Y2�ÂL��o�d�e
"P��lRg�!`BqU���$,���}��'S&��$岷22��ȅw��Е[�n��#c�W-��%Ґ#T|�ͦw�~��ϓڬ���a��+�:P��4f����]sub��-��lX����5��	����!�(0�v��8j�X���L�:S���d�.�#�/Pi�Q�.�0w3�7���p��EPy�xݯ�A���x�Z��ϕ07<�U���47�QK�t��3(:_���al�_�J��,�Q��9��e��U@�M ���F@|��Qw�86���t�ӂS��*�D�z�����v�k;5q����U��J�M�d�<��` �>H!C�<��1Ԭ�a1J�G��>6b�/a6\�9�AC�:����5k{7Eg��]�֚K�MH��|��;�qo�� �̐2E�.y�K3}o��P)�G��dDfU����F���b�ԌP�bY\Y�@�VIo0?�i�s`݅[�{�����w�V?@��J�7�|��AG/05��`w�� ���0Vt]���E�i�T�.�%���_��F��4)������>Nr�a��h���e�=��dEg5Z��k����V����e�2�")��E����4I�m�~�>��a���t���&�?E�G��H��:�S����hg�1�˵0tj��iC�������i�aM3������*���?� �s�eB3�]X|.��8+��듅�P'?�Hǩp�6�o�byx�kP�
-}l���WG�D)juԒ�'lf�p��y��"X�a������ݞ�jN#��� �ㄲ�y�~�r��Rj��3�i9�8����U_�2:m�F��W��������܉N����o�@&bjf&�S�M��E�![,�Z��3Sjؘ�l֣��a7��S�?����L'JFB	�0��<��&E����xˆ�.d�1�#�l���
�E�*B���sp֠EƵ�S�x�pC����b%�
���(&��4
�EBGQ�Q�AI|��-�#{l���v?�"R�4ve]|�Z�Gda�v'�	��٫*�����nnM��]��cS�z}�*p�cHe�/
\C�ѨY+����#*n�öw^��Bm'ss�ֶ�s��1Y+VM�U�j�^���h7>M�����?�>٬UV�Bl 	DkW.\`=}I�!N⬴�g�-٩�3q�;��h-���������5.��4��l�w��@��ilD�sH�y��;��鎾=_�n�g�����Rc�'�N�}��I���G�������"
<���:�7)
QvGbC)�+���'0
�ŷa�H�Y��S��=0��K�_���g�u����Β�"���(���'n>�v��L�41��yv�n�c�C� �z��I� �ra���,�c���;��ˀ��ğ�̐��'&����8"�r��T:Gv�^�T1��/�mI���H���C˩ރ�N�s�KYY|��7�jjI��+���E)���U�|i����B�=����.._I���W���s�=}������Qy�`GVU�*�!���t-0��.�76����se����@g�#�~;Խ��`Zk\�~�4K���H�φ�̜v��D�uA�/�З�����j�W��]<�~p*th}/�還O>+�az�}f���,�}�|�Kg���v��ja�XD�F���`Tr\�y3	�Xy�+����Z������I���u�#�.��2nG��;5