XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b�E=v3����(U7��bl�dri���a�2(_/�;sӢj���W���;��ٍ��:D'P��B����1d�����qz�bv=!�z�h�7c�a}1Oxo�(Nn/>(K��u����erר0��őO Y+^��LЏ�G]����Qk䲔a7�4�m?�	��#�η�((;?�J�YK�-j��ֻD*U�0��3%����!gTU-���0`��A+Z��c���v��e��:�e�N&1 ��ݫFˆ�>��r���]����>�oW߇�+�W�[�D��ӇR+\��Rm�)��C��v�?Ӫ�C�;�D7Y��,t��wP�r���6��z5�)6o����W�����������^%`��`
�1^���b.,���C�	�}%�id���'��h(ʀ>F)�>�i8*�I���1�lG�"6�y�3� J�u�=� �G$��[+ֺZd�>�2�m����a���p���d�;s��O��֒�N�3�)Q�Sw��#o��ZP���"cBDet|�-/r�Mvbg���=w��`�]�	����YA_�n�F�]2¯���D���²����гV4�����Y��yqj�ňT�n�߆��|��Ծ��-���̟�EeKѾ"�<ɼq�(:Ű��V�O�/�9z�)�eN�+
h:U8��kY�J��c��B7�x��F�@�`�}��&���=j� �G�=�@�{�Y�gH��m9�$��n=�
i���UCڦ�T�:JA4��AQ�>�\%қ/XlxVHYEB    5224    1740�о��%@qy7�7�6偤{�5�w��n�mF��t�����-�[t�iL4~A�
tQ|z6Jw��CK��Z��tۯlت��'�q+*$#�\�	tͿ�e>�Ec�i5ob�cfPHҭ/�i�L1FId�B.˙��W�����E�Βm��d�d��(_c��u3]����{�H�HEaU9�c�Ck��w��(�h�l}fk�ی�=C�4��h?�K��48SH���B�݊��}�0�-ΞlZ��0�C>�~HJ���t�7	't�o���B���(ò�q�*�ڎ�V��/�e�B[L�'�?"�E���a�q]������;g�a�m��w�5^>f��c�Sx���_odӂ� L�C�h�� .x�Z���7�_���a��x.y�u���%>1�J�yQߵ�hEjY�j$2����6<�޶�C�=�N� 4Z
8?�y��Wj�c�#��9Ԗ&r���RYN�2�4���/�ٙ��L���y؆@�|���(X71��M�\;\BT�!zn������e�H��LK]-@L�B����`��ܣ���ˤd����k>��T��:���H(�;��Y�xDcT�L���"|�4��I�Ӛ�h)��?��A�P�d�A=�u�RU7��A�:�g�pu$W��l=�� d���32d�'�=T"��.�Uuƪp���Eg��&���0���Wܔ.���Ã:�����w:��6eď��$�5�~E����=�	V����k�eˎ�z7��f;8�nQ*]Ŏ�dY��2z��A���y���F`գx�
_��\E�1���?���W}���_&^�L��E�� ��� ��v����y�i?����S��]�]�7C� �� ծK�Q9� `����B����< ^��r�|Ej��w �����B�v���9�R��|.x�4y�Q̻��nТY����6��@z�(���/���	mF|�t�7���B��"S�j�m��!��C���C0�Ȇvf�I�}�W���}:';I�T+|��eUd�H�N����n�so��w�	x.{������k�fm��H/ ϻw_s������	` ����Xe�9�j�V��>\��:�����k		P"]k�Q@�)��p���6���#���:��p�R;F�������R�;:��+%�^.%�,U?�����6�>���P�����$�o -���;�>�_����:
�19k�	�C|��O|���b����l�,f����'����gIE�fZ��S��%e�Bыx�׫��C1���7���r:J �3n�+-�@��=�G�MP���}K�2rj���r��.�}�];���Е]��J/!�Ü��u�|�*Y�w+����1#�V��)Tg���O���|LW���Ы��
֣�!�!fB����V���E�E��;7U�)�/և$����I/���K��b�L';��
}���A�I�J�})(�E*���k���D�;zz(�}YG}�ϻ��Z��FCH"1�TV2��o�0G7�7qi@��ŵ�_��w)kP�������	]�(�c\�
Pm��y�S2�.�b�(O�gP�<�N_�3�i��Ms���%�8��H��\"R3�V�kM'�2�jU��h#�[�iAMʛj$_�*�U#���Y����Fz� ̺*�������e�S��M�U�kO2�'y<?���
<�A����&������GEA��rP���k�P�Щ$$.�q�18x��kf�;�]k��`� *O��oV�.#�p���1�3�w"`�Ԇ�x�e8�%�X$q�;1'��R�p�,N�BW-Տ�J��'4�H"(�DL�E���id�Pax�`�����儲�bū{1���*�Q�4�����ζv��,~mᔵ��R�0�M0l�[r:�e{~�҆PbBf|�k�܆�)F�S��D &���]�ɧ-/���{ۅ�GM��Ck��>3�����o*�$�;�����!�9n���Sg�G�S��<��s6 �ӄ��N��b�ݚLR��$�:l�.��P��v�R��!g��k⮚Ғ�̂����mE(�3��3C�zY|hL#m�Z�W�FFb��܂��8h�vz�Ua+5E�*�~@m@2�)�yD3M:�!�
gn��v剏���r;�d+����O���Ż� �;��𷏙?E�y+����4E�9��C�$��a��6�Ȧ��P����Y�R�L?��L�In�%�x��*����n�NnP�1�Z-�*Z�Cgr"���:s�MF�j>�����c<�����z�Ɍ���)�3��c�S)6�X1=�"?��A�~��9*;a�d%?�����Ȑ?)�8����ݣ��t�R���eyj�F�^��tx��;�(��I�Aw������6�K����C��@ON�����(����Ln�X�+��(6?�*H����/~�S
�e�@���ع�1)��$���2���~��
E�Y�%�ݫH��3���z�Oo��7�~z	�%W���1��fXs��w�#)���$��@� Yn�0�:��P�#����ɴd��)u-�����%���+Z1�_�����Y���X�$�E�p�Pɉe�"])_/'RصV�[�����9z�.d?���+ک���t�ε>�S#�s�-�8l��}�>F�ڢ��%{ha��3������D1��3�7ZR14�m�(��}�HGn'\�N���q�Ѕ ͣ[��Ӌ��^�?'	�����SP->��t`7�[vz�;-N������I��VlQ��w�����^x���r�~�/�H���i\㦇 Rx������s�D�w~������������>�%�������\U\[ky����^��T=l���Kv���j�|z��qڡQ�?��Vx���Z(��D�p��1��hʎ��$��18L�{?�XO'�h7U/Q.\��²T��[m%+N-D�B��P���C��ȳ���≮��I�F��-�6�-��C���si��=Xp
W^�&"���V;��y�eGwc�T6_�:߬m���|�j[� P�j�����I��(�k8��dkQx���q�oE�n`VJ�D8^R�KE=���H��U���%����a&�|�>� �?�:���ݞq�͊�m1��+X+h��}�������C����2|��7�b(*s9Z�O���R2єv~��>?���ͧ�B�Y\L{���s�"3�/36^��s�y0S���;��(�w�׸��>�ŗxŗ��iչ�X~_�g��ejork˂sFBl�t�=��Y}�
��!�{�wȋ��Q�l.�Y���%�h���GL��o�VÛ�M�,B4<(r(Fd!�	*Ϳ��sd��7�ʫ�M4S�X�ދ>�prs��N��ؽgָ1=̞o��2$�ʭ9�HN�詏�F�\�@��ej.Dn\f�BU�?9U:�����R�Kf���u��:P�S(Jc��m��bs�$��O�.�c����?{�|����Q'�����%FU��X��=�ǳ���e���T��{�!����(FX��85��ڎ
z��`�u��s1���_��,@G��3�L�1L�Ǭ"d������l	���E.����z3f3�+�N?��A ��VY�W@{j�(A�:hJ��+�Ҧ��})1�¨P��5~
�៤�$(�F���\��Ȱ�>�̉He�5�J�@��͓�h���Ot��^����.�5q��8�Fa�ak�'�zm�|`2��T�h\諵@PC��-�/n��}�@��v �I6n�>�I�D� E0Z���~J��6tc;eW���k��+\�X�w��2�FX��ҿ���8�9 ��m��0�,��b���!Ȁ@@�ֶՅS�	�����G�s:k��yY6]P�5�4؊�^y�_9��G6�^�}C��t����2��QoC�I>�,���7���%�p��#�`4-���)H�˵��1`GI��1l�cO�Q��}�#��<����20��~%"Ԫ
�!���,&+[��}���j^�4�fx�ɶ~��Ƴ�DkS�C~AUw�x�������/_��@�t�>\���V6�)�P�':�T�KJct<����(�m�y��˕���+���R͸6�1�U�����%�8�,0�6�#+;h$U���|L����fzH�����f�ھ���"��y4IR#f���l ��v	n\�W>6;$v@QQV��p���=���y��E,��	AL��l[�;���Ьzz������׊�j6��l6^l<3�q����C�g%�9����9�-���.�H�ĿA����)y���^ q<�ݜ��F���B��H~Μ�E��E�M���kڛە���Z��U������F��ۨ�<���,S2�b���
+4v�<��T�r�<�Gy�ä��rxO4��~Pv�,�0Ϗ�1=�$H6�"4Py�؊�$���̻��<�P�ƞ��e+�ʱ��w�Z�Ύ{2T"���?�ss�e>I�xq�DU̸z��~�0�����'���Ό{��-���݆�NbuHΨ�4�m�w�;���t�� �\K�MH>�~�1;�oֱ�M߅1�z��
�VN[����ʯ{��%3�r�}��-�ok�Y%���q&�����.O�G"�0���Nm��wX��PH���Giݝ�,��������\�23x'������>٤����Խ���<qzzN���I�U@�W��=!U�%����(=,�&�!�ؕ�Q^���vW-:�DBP�d��Q~a��b��]�}�6N�6.GZQiڱ%�Ta]�*��"�K���&�%V����Mҋ���A"�8��^/~��C��ٵ��m�|/_�liw�
n�O�MB(�V)�$�TM�d���J�~y�������kI7��� ��MYU��	��\��7�Y�'�A��t}�Â)�͒;����M���ٛ���q�se���EwS\N��*�S�<��=�k�� �^�M��y�p�Q��_�ȏ�%�|XT��*x��,�罾��]6�S���U���,�O4k��<��D��D�B�=r���t]�^:c�K�J���&�mlFs%�-��	era�Tk+^UtSүwd�oD�d��`��Do[[5�`^�H~�QM�/�����t������pELl�`�0��1���.pikKAU�a�l!�XϺ����8�.^�~^��W�ŵu��*�$�v�\�s`Ũ|���&��U��˖�ؼ�I��iK���@���)�#k 6����� ˈ/��?��V���w3~�P��i3̩��j�Q61�Х��m�-#�<����>+7����T:�D�w�]&��YK�^��Y�;�t�1!i�Q���MG��ލ�T�M���)���e�4�;/\�=�!��;VI08�y��
��������f5/�&��xe=�F���!�,������E=�?\7/�+TS�x�L�S��'��f��za��_L1���.ߧi���׸��2��I�jWg�j������fؤ3	<���5�N*cό6��ȖR�ϳO�Ȼ����(�%"�ce�Xs]��3ە6���.��]�#h�l��TO���i��f5�Sҕ!��Y�IA��N�ep���p#���y4*|rʭr|�KE&�f��?i�dژ�kW�
��w��AA*���7���l1����\o�vE�n-��w�.�:*4����7��x���騰C�@��C�wB�Np��T"i�Tr�ݰ#�?�شm=\�;7Hge0��u~�\�C�^ç��sY��1��DӋ���6w�F��D#"3�?�]i 	P���^�B�� ��vw�$��x��IBG���M[�MDS=���	ȇ�|�ꙙ�ό]lQS\IW� ���֡B����F�f�