XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���B2h��x0�͑Ab΅rRS;>���Ȏ��"�e�'�o�?��_#� r�]�QUPz�R��ȍ��[<�۝k�������
R��w_L�b���E(*��7*���cv�q7��ƕ����̔��%�B1��k�D#���^����� ;���ڽN��i�;���H�ٕ���Rp�c�и��fRwM8�U��,�(���:�p�K��5�$��1�!����#��V�jl5(�M`2�ɭ�mp���o��2��6P�:���[�{�K�T��i�
�˓csU���O�,o��f�X�1�_r�J��
o=M�i7�w`՜Ao�Aa�K�{Y��hv�cvԞ~�e١$��%�̡S_�1u=��[y]����gh��.��r�I���.G����]�h�f}N�����G�l�4�&��dt�1u4Ұ.�^�}��k�Op5��q`�CL���{M�������<?cM8w\������sʊ��,m��h?�f#ߕ6�OL��&k9�v��}�7pd!`�37i��<B���aG���s��N�ۍ�dg��{�~�������iP�N5��"��O�M��k����Oe����j�����h��R�
����o�	���t�+T6�c?hg��`+H��t�n8D�5�̊�n!dZ��`����������ړc	��l�������{3.�bx��N%�Z���q�
��55�̒6{P��*�7w��ڀ�[q��m���a�􍊈�Y����c�/�o!��gXBXlxVHYEB    2326     980���m���7^��I��:����2�I @����7�H^yxS�h&�|���h�T�].WJ�nn�sp��)S ?t�=�ly g.��f�IR3\���������	R�9�S��rs����/�*�.��K�#��]:6UAQ�h�ٹ(
�_�m$� pu�/_�XWP|R��mh��v�zZ��L���u��c�?��73�X(���#���:���-G!m���S|W�t�
�N�Y'�,�B�E5nI�ւVj��b����AOmJ-��2�K��v=�D��p�Hʌ�3\c�s"I$Oq�6*��K�XP���b�&�8���#�CN�;j���*���TcEh*G���AG?_�i�\���= C�
pw��rd�"�W,�2"�F��;�O��k�ل���c*~v^��=�����a�3[N3�rZ��F<N'ے ��ѳ��v)�(�=0$��_���R�p��|���_���B��J����!�|�y��	�UD�_���>�c���� �xR��D�$��Ҭ�[2m�yTW	Ê����[�������`Q ;���o��iT(g_B4��R��/f��� �T.�-����\�Q�w�Ѫ$ֱ�����/b�1�r��o��4�7p�_��<W�T�@Q&1S��4�N+�@"��41���8��}3k�^�%�a����SPsZ�ě.�7C �@�@�ڰѻ�*��z�U[��/,4�P�I�6`/5fe'�iy��˔�J�^��KV���]�0Gdc߁-�͌�����%o��g�[���?1Q����s��\���^�l�4d���L*�_Z�|���qO}E�Zܘ@]u�g��A24c��WjTf؟,��aQN[�xu+r���>�1Nx��"n�4l]�4~B��=h9ƛ���8a�K�IX6d<����o]ɋ�P^P$���ρĶ�Z�[��܉#����V�����zr���yƜj�tM\�e����l�Z�u�w�=F�v�+�
���M{�b�+Oz�Gw����r�~�Eb��v`���:.&[��S%j�F��c�S#*��y�a���,����ɿi�-Q�|Is���K��u�����8����J7yWӠ1�{��9m��`*���uLkF��2ط�z�.�Q��K1�Ӝ*��E�tԞ�}Ơ��i���̯�<(�ݔ-|��]q��n�'Bp�o�8�>����c�3��-���W�N�4�m߉��A�&�� ���v����v����H��+��߮��e��c�;dg��纡��XK�:�GFS��pV��!��)���S�i	,OͰ���2D�tN����7 V��R W��������e(��[&-� �.Pt�G,W�`�7'�\6W��3L��
.�;I�d�q���W�$���JL�X8����A]VO�)Z��'b�~?�ޤ�e��J�����9i����Vڕ�@K}i��7�}��g����:�?I������d�Pa����r�̵1p��>�t�MrE�@����ǻx�v=0�B#=Bi�S��'ӳ�TxTJ"V��0I�� Qq�W��~/f݉�K	��\�����As�`��v���w�����V��$.)7+OZ���f��Ո�a�c`�ُݱ=1��j�$����l�~���.�c�2۪��I������m�a��V2l�B�����Պ��QXo\_*���w������f}(�{�����m&�w#��_8$�ef[S�'P��]��~J��L�	��>��#��/�s@��o]%�X0qJ��.���g�-N��2����x��Dߍ�I�s];�. ���ua}�ϴ�jl9Oo�a��~G�i~���LSwB��O%�fѣTC}܍�G�����y�;{��_z�\�:�2����ޟ+X�I�=�/��~a� 3�� =�Wl��x�a���H����F��6o�%�i�~�%��:��;�y*Ґ_>g�Ɋf�4�]�/�S�g��!8��4�x�G�.4~�I�/��WP�֔*>"�1��Ќ F�G�)�Ã(�D�#�-_��%ҧ�(8�ni�����2���GV��Xf�C�� ��������������э�����X�u&/�Rf|�����Q����Z�gt�ǘ�*;�����\R�>��Fh������0E`󬅙���T-�.NY�iQ��������>t3%�Kםǒ�ߏm*�i�8��TF�h�*ug��D�`L��UJ��5��O�,f�>TA�>����ȞD	v�mOEe�|��Z�,j�K��e�k$,o��d�ۊ���� ����z�����ma{�i��1��0Y���hL�!�>\K���D�d���!�CM.�nkq-�	v��n��l����ʪ�|�G�>�lۢ��8Y�6�#�淜��������x