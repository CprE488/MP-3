XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ǅ� ����g/�~����y�ہR�ٖ1�B3�k�?m<�@m%�%�	�@o.�r�����]$�m���`�Th&?6DR���	�=؀$��a�CoFx�kЬ���k�6�X�{)���/Y�#h`��R�.�_p_�;�йn|L�0�r%ڙ4�6nKP��˪8$�Og�.�FWzk[Mp8�ĝ�oD5�����"�O��� ���� F�]�����Vp��l�\�N��E��qJ���Rx~b��:שe�M	��R(3&����� 2���

VR"  �\K����P�k�Y6�y7#���2~x���JX�%(��t+�t���ӑD�v&U��#����>��C�$vy�p*�u�	.��a{¡�o�(b���4)���+�4�e`2y�{�1őn����U{�T��c�KA��`/�"�^�;O�{��yj��[tYӽ�Y$0}�7J��q"���W�i�h��؟��#�Jj�.lĄ&	�:��ǦrZ�^ �	v8�_��^��%ƿAυ6)�*x:~_��V%���#���Ջ�����MD�EF�=��:GPPklwp~���k�D�y�V�]�s�T�J�"��\�eNaxv�JF����E�:R�h���[�}�UV`���j.f#���}k��9mG�\3��D�D�ȟ!������2/@*�	,<�Na�.)yX����y;=��˒�v��X�B� ���_��z�Ӎ�L~�v^��nP� O6�4�11�^ѥXlxVHYEB    1e3a     a20���>/�M)�*������4�(�Eiݻ�g��Z�߅�I{�q���Q d�C�]7VK��'.�:Y�5�� ����ۣ�;_X ��)>��d�Kv��J�Q� 5��?�k��I�,�SdfeЫ��4�k�Lӌ�+23~�o(��̚"�v��G ��\jO{
2 긼�ZQD�>��E���-ϳ������&��O�l:ε���J���W}o��̡�G��*�(L�4U�>_��X�W�g�����"����S�,)]*ώV������C�=)e�* �H�,����U���m�j�!���9]�H9����:l��I.0�� �a��0���}|����A|�!4H��/��y�J~L�iu�W-����AP����;3�Y5�r`R9�\)5�K��Љd/N+�����M�1����;�Ї*FE��s̰�@
c\�M���+�<_�)��j�rl�E��"(�_�c7�x8���8�_XI2P�����2�������(�%ׄ{a��0�m���S����ə/�R{)�������"�嫦>=�t���<�����΅!��y�����Α��]W�Ս��N�e:ٻ����N���Z�~������w�F4�]�q���2?d��$X��qXa߈&�fw�D�wÆ\���^��a�R�L ��/~��煨qhN��BՓϐ?��y�l�_��'(�$el�C�����_��c.�i�2뼴F� �͵�S\�O�)o@"����?"�k"悤C�/��'.�}7�E�չ�#�)��\A�����w��=v�Y��}5*�fϺ���,��Ӊ�~J[�N,V��A����_ݱ��#�V���j�� ��)E�@"`3E��/i����2x�f���F��@��Q.Ɯkx����ª�>�l���H$>�F|_Y��`h����fJ*C�rUG#�%cE����ƥj{Sۄ6����Q�����Iw\����W۷�uv��Q��d��;���c����>�����M�rʄ���D�6�̓����9�$��4}Єx��+�|�n���E����DI��J�n�=��t����p���K,fT3w�<IR���o��?�Nvl��j��y�ыR0��j��_�|��
��%W��1������Q��;�	b2$�7�]��iy�*��p��2��Ne��e���&�h��T�c(��V�b���hr�
�ռ���B��į�0��G,vA������G��łM]/$�s�)u�����pya��,��v80�X_��˾Ԍܯ���9�d���;7�؊�3����YL5�������:(�
����x�8h��y7�j��33w����ݾP�<:+{�"�e�I��(�9��9�+����H����OT������R\}q/`��W=�P̀7�<�.I�q\]�ڤK�N�ѕ����]�u�Mu|�}B��o�C��5�Q2��8�z�B������j���� H�2?���4���c�"�f�KBM�Bф����݀t����"`%<=�����Ip�_e��	f�D�V�YІ]�d�t8�,汈���7��M��T�cU�^�ˢF���H"�})q��jC��B��.���MT���2[ �$��0�����#;����+p3�읿�p��S��C(l�����rgY�{�O����W�olɗ�>b�ر�����}��d��Ihh�j!��B���+�{�~L
�||tO�N�_������ל��à��.���l�2ש�U�Ź=�@J>��j��i��➚A4x$�7}�ڍa8r�<eox~���l[���/X)�׏���� F��Ⱦ�a&��:^o\�mϨ΃�#�&��]���&/���W�o�i7��!J���B��ƴ��V�@T�oy�Ve�1�!�����i�J�p�6��{�Lσ� f�X6S<��<�r§����_Ǡ���Sv��)���^�;�����Z��`J<���̣:�V�t~��1����F�\��o��$��h��?���u�P҆���1(/{��|�*,��9�k<Cw�9b�2 2_[�)�[�m����P�U@̪��x���14��bP��WW��N[��x�BLd*�\��t�Tb�Y�(�Мn'���e��!�"8�jRgd�o,6;	<Ѳ��J>��8�sQ:��~jY�Ң����c��e:�K������,�l������ߘ�4*y&r��g�a\�b���e��_'ɶ/h�G�T����\&4T�C=���x��A���˼d�ce�{��{���z�H��WQ(�ű�{ e�����c7[�����햫S����������v.�t���d:��Eu�R �t\��K�ߨ�P^��#r�Pнv���o�52��@7�_j��qP��q�Q�Xp���8�P�Ja��}$�e���̘q���,�;
V
�(U?��0(�C�xft��Ig{� �5��z� Np�F��O.����4�;C������'�1k��$�پs"=�V2���A�O�;r(�w�)�ܚ��3