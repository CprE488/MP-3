XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������ XH���J���<Dm�p�NZ@9���+|�b���63蜦��K=T�N�R�kZ�6'f���N�[��l��L�r�T H�7��<�_9H��6w��;�!�X��w��N5H����=c�:�)Ԫ��_{H��N�y��.SlK�rW�JN�Y"�7��"3��B5,F�]���2T	-�L��� �t�tz�.INJ
Pc����Y϶ .��� ^X���dA�r�Yp{6&޳��#�T�� ��̟���w�c�o���]5��������ɍFǤ��M=eN6��YWIèx��5 �=E�tK���l�w�MuAD��-4鋍�Z2��������b�=_��
��U=��
��K�@�J� �\"���s�PmǙB���,�������ѿ/ڗCM�J\��I� �^�ztt9��[��s�2��Z1�纟���Gy!@v���hi�,�}<�eصk�[j$Vk	�"橺��=�}Vͬ�n@u��cDd<1]?�6�7N��Vmֹ-��fh��px�Oi0�ޞS�bh�`�X �8caYv~���Q�iTh,����S?9�q�$f��M�wf�nq�Ej�i�e�������m�j!��_����=��qJ�f/�h����&��ҷ��S�"V�����:5�nV?/��[��s���1>ԪkLG!AJ��j�п)���܅l~�FR��@�I�J��]{'G���LHh2Wb�eݐn�2�:�.��=����ߒXlxVHYEB    fa00    26e0J�z��da	c���t�/�����#�L�B_�0,���Z�N��cT[��eh��'�1�'��V��x)8ug�Hk��d�v7^ן. �s4��t�J���
�\ͼ�0�Y���\�N-˔���F3�o���4*)��v�y{�E8w`�vl���yn�Du��Ѡq��M����at:`@��3�q`WU�f�/j>�"M�tMv�qg<���Fv�vb�,M%��0�7�	��$<cX@�4 qJI�P�:T�Ƚ{?f�e\��//�u.��6;�2-�1攪��>��Fp�ɵ�#$7$ְu�_��8�>�bl�O�'�4	�ڜ�~Л��g ��|7��yѽX��L��'@q�%Ȗ��a�w���l���Y|-� �"^������^�H�U:�L�d[���_̏��
�T���4q�����P�H-Wб-yDn��W E!���D��U���h�*�[q�B��V������P�d9L1ؐ�LEUUa��F�!��*��T�I�\n\�U��1P1L��h{i9����q�ܖ@��1x�^B��w$�Q%�o�;AY�]dN&�'��K/�}�-�C��GmP��r0��	R�h�R�WM��}i5')�Mq�kH�������?L��zL\)י	H���	��l�G+q��LO��9�5~�9��S��@� :M�(p��w� {o��·��g���c�A��! b��\!JW +��U�8���v�XQ�0]8��뛋���\�`X������0F���@἟,=U
��r)	�<�߄>�����c
�@$��M)�:�@�4�4��@�霾�?!6���Xw̛�䐗�ƞmB��	r��(U��{R�����˚��sւ�^������6�|4Y��[ ��+*k��G����\��J����@�)�� )�<ᧀ��-�AF�m�FϜ�&���E ��'��aw	�M|~��fO�K�"����X�+�!�c�����;��DZL��껣vI$v��ӃP��l�$���.�f���5��-)s���R���n�@�eJ�p��b�~�<�>��j��O:��A҂�����.&g���RE뙽��u���*+ϑ���y��}��F��;��&g�懮
-�A�����n|���_�L:I���Qȴ����W�6+���y+x���&��.
GҞj�n��n'x1�*���Y��Ԁ�c*���c��0����X���;��S�dzlHe��9f2���I2��D�b��Ȅ23�{g��q_�
�$}>�ܗ�3�>
�ZQܒ5�DI
5Oې�]��[$C�
��h	Z�$�K�Vt��g��֊�*sp���v��C�6�*a�+���¬=I�uh:>����X��&ї
PR�3|�����*2�>6s���}@�$����Y�_|.�_��y�r=�/�1Z� ��$�<(�D��~�g��:y@�r�;}�D\��ಈ-{gՖ]����S;ʟ�b�g�v��jO��Ç�bD�+�tz���n�ߞ�x��כ3N��<TE̡�Z`��qu5�J���hV��?�&�6ihP*��L�5�R��ɂ8-��K����C��Y��gy�)�����f)��;�K��w���4�I��zٿؑN����.��|0˩+k�ì�9K��@��	�%���[��?>4�h��}�����p3�k��������_�G7�j_M���@�ٌJ-.��˕$N,V51��^�ć7��i|/��Q��XkT����K�yvr�+��ai'��;�\���6����'��T�;�|�Xn�M���t�{��7A_U����:M��j�_��|8Mͷ�/>�ǬΪ�$���� ���ɕ��F�)L|L��Ge�j��0&-1�
�������x��Ĺi	�$3�?V��IN�'Х��[q��(���BA�4<�4u��9���9�f��)��M\h�'���s]V�U.O�׹TfS
�m�F4;j�.�_�����m6UB0.�9��ʿvR[`���s3�9��5�������q+:�qN{�7t����'��)�����Y�Uk;�y�k$>f��A���x����ky�~?��rX���\�K�Ցx!�CK�s��i&��(g�#Et���Z$\iI�z��'���h���zTG^�5��rC��$h�kK����OPV;wH=���w�3�s.������|��L�u����!}��SE�#��zP/S�]3	����ʓ�y!;J�y��kukя�n;�h�����û��G箛�!7�������Fq��ы� ��t0��f��Hb!�/	��ĥ ������$�޻g�h\���w����M�D�:�g�]��g���Q��iTil��Em�;��ȍL��0�m��}�������a�?}>�8RR�eÌ�^~�[nU��+;X����g�R�e�4�9�2��4�����/�ީ�.�ޥ�.��d�i$p�Srp���:�߷�ȁ�h����&�c��r�|P�h�Vm�Y�v�[A�KzK!j��)ᤵ��8+�ޟh���3A�)�nj�Uţ�	I�cO�X���|1	~�?�" u;�I%^'�]�~;�Ԗ������MǝS�X���x.�*b i醑(� ̥��ᅚ�!ӕdqXlLՇ:h#�f�4���6�ɧ�Ē?�2�eB�~��V���}�TjZ��tapK��6�����ٻB+��jj�b��`n�xմBAf�N���>m5�;��çJ��]�,�L�hw��+&��i0� ċ������ymj�R(�h�CL�,����V��o��q1[�&���e]���IZ�n�&����a�(`�Gmj��5��֒4��0�� ��?)�g#��s�˄)Ѷq��e�������l����AZ]K�e� uD��8q�B֕�ub�Ǵ�/��c���-����^W�+0_	�hi@�f�]��!����]]�P,�g�D~0��rO�9��F�Ƴ�-��v$.��	�����F=/˻��,� �g��OR5��Ǵ�D���(�
���w������0
�$��H�����=�y�^:&����2���}�m8#&q=s�Ь���s�n��Fc�j��4~�w}�AVNAF&ԃ[D�r%ْ?��e�,��j��G�T��y���D�ZES����5W�⠓3�� �z�P�P� �>'3�VlDM]{���	�o�e����,���e��+�d������%�#Ey�WC��^��[�����n��PBy�+i����/F''{�����n�6�nS��ل���Ӣw'�`HƋ,�jΧy��5��lV.�goKl �G��{�4*��DL����/����o��o_B�;0�;�a�O�v?R\�Wr!���U����KI*��I�h^�١䩆X=�NU�zX�M���mQ�
5j�ky�q�o��-T�ꠝH�YFeԞd����G.�;zD�35�|{K��*���̌���b�XC���d�{~Y�)���1�C��˒���Ӎ��XR���y��Ǒ�[}���=
(�<�<�O�u:��	_��@�����]%������8�o�B�+7�o�A}�4<��(,J�ԕ|�'��i�6��x�ۣz���ɉ��?�Qp�;���4CE^��yUy��UOBQ��\T_�$���(p�-F��O�0�2)��[��S"��I���]х�������N�8��R�=�`>Z���Ggz�Z�k�hS^�Y�	6tQ�/���p�g�4�'zY���9� �NAQݥ�j�+���`Ӥ�r��~"���9ڭ��;���o�͉C��+*�aG�·�@(�tB�Z�V]�!5K�� �=���ொld��n
����uT#�a�D;O��MI+sU�"D�?Ȓ@i?����:U��\m"�Ձ����FC���`6�4`7���?B��ՎQ��L����i����� �[e7��?8������21���3��Z~/-c������>�`�� �~N���P�X��0P�03���^9��_ȣ�ƆGFm���#gɋ#��Pg��Ӕ��oY�Y��-�W��Q�8%P��1 �_,P˴��xpr��1~�!��]��UT�D<�~�������Q���<�R�R�������Uz�xC��,�Cd�m�Jl�nX5��@J�d�y[�j����]�K�Ɗ������_�k>��M��Vn����X?G={��ART�pλqzF�̨I�����S11m&� �y��Sylna]u�.z�5K�)T+���t�A�*"XCu(ۋ�^6U����m����S/b[������a��f���6�K>r��H���7�
�B��VA�GkR!���T��5��,��=]뱛���s�$�i�z^� ����\���F���^�+0Lj�.V�V��Nl"r>=���#��J$]v�r�))Kh{d8�`c=s� gTV�"y� @��H�l$EŪ"�x���O),Kf�BE:�ѻ\�����ěoY��㡚�E�*f)�e��6�L�.�����Txհ���/-4� D֓ؽ�7h$}.7�$Vjk�3�1L�:?^�>�#
l+��]����l��J9�R0򨓢�Г�L Cf�����R��ceP>����] �O}��שV\���C�r�i�B(C1�:?�2��eWX��}L��Π9{�ev���ĉrYԧ�+U�9�2�Y��n�xX���]sh�0�?���� y,�v�ز0]�چX��U�]KM�S��T�g���L����r�?ўQ+�*I�E�_@o<��)H�6|�7ZOc��D��r�AҖɰn�S�0
H'X \rc�r���;�K�Ե<Jٞ�9�wj����������@;m�������@�9���:PY��A*�����LB��O�Uw&�}ۘ�1�gs��I�,��?k�L�YO=%�B�M؁��ې��S�I���b
��C��th�"�`�3�=���#2���Ӓ&+�3 ��M����љDʴ�~ P���|p�y���q�⍊8S�a�TshBNC����	w2��S�$GP���%�p�X�{�]�if�Ջ~��JW���B�w���g���|���=n��YdB�I�5�]���B¨���0e%AE��e3�|���U�z���o:�?b#���S,ƭ�d�^9'��9��pZ"��7f5��u��+E��C�l��OW' �/��������GO�<P֥	9۲Z��>���oBȄN8�YVb'�j^]�B�Y̜4`�/.x���8;~��^xXam	T��؂��>�t4ԡ}�4��`-
Gp/�L�K����>�8�ΤY�G!,vy�+?��L��=��אCp!l����%͍����蒹<ZL፝*1,GO��,��ppO5��_��P{�rX�T�&��_L�T)���W����w�1S�a8�XģwBq5͍w%�D�Ui�NI��A��|H詺�:�������|��6T�Ort���隈���ƶô��>����.u)��X��G?B��s����U�9�=σ�i�ȵi.I���b궺B�CZ���=����x�}`vd�3����!�2]�Q���-���n��/7�����(��l�كP���%��-�����5J��4���|�~�.8�
�)P�SkG?;Jd2�dϭO�>I>;m���2�2�g���uR��h�CihM����c��[۞#�I?.��41_�KK����������x��&<j�J��i�DI>�����QV4� k�!B0n�R�&Wo?��>��~$�@:S f���D@$/��,������������2�[�of�����B�+A������+۪��;�A�$�Yiz-T(��!;W	�荄}u�M���\���M��E�9�I�{�lp��ݍZX ݗ ��I)ᥳ&�Q������&����0�l�.+�ˋ���8�"�d�Y�dm�D�&�O_� Y�}Bn�7�S��~�I�8&6�>��S���N��*r�O3�88�T���g�j�k�@���i�NUܮ�x�~�(�-�F|?OX�(|�$@�<RZ�=佹 �,
�C��d?/�P�8��H؇�M�#}�8fQ�(�6�������^�8�&�x�ӋѦ���i���&~����H�hs��0F��AU��hu)��}�4���1���.A��/DrX���;˗��m��#/�¨�k$T�8��S�(���������&�9��@�Hpa�0�b���IV.-X\vJ%�?�ά����=o���:L�������z��Xuo�5К�x�.��H��W3m������gYL��P�W9�U>�)�2l�?�=�������廉ޫ��qS���-c�����@Z-jၖ�?e�7Rm�W���HdkٞU!��N��7Ȝ@�4��UC�[�� Lh燢*�7*���.��6Hw�V!�F��\��d�a[զ�1�@c�DU�;���;��i�zF�B�V���!)��l�b/�����"�,���5	�,4cl�D�h�5�Xň ��ߚ��l���N��X��BX/�A�:�.6�g�>��Zh�kM�c�ۚ&u/{�#$O�j�6y�}l��AS.���:���#�P������W_�{���C�g����e�~� Ԓ��x��m�1Ǿ�F6��	�&��]���C%�i���%���.��F�:�$e�W��/�IH� ����K�	ZՑ�Td��!`��Ȳ�s��p��/쨣�:�h�Z�ߡd�L�S.����%�s�-���ec}�Ž���*��q)a��� �nu�Dݟ$�,�:z�9�!O�T�"N��)�u/<��'��М`�tw�0��-�/�^N��p���B3���y�j��̦�&�(x��Im��
=W��:���O"7bq%���Z�2�r%�9#�!$�K���Ag��V7]����s:-Vg�����|=Ԫ���0��H�k8R��x�9^�I��5����r�>�
��3��~�r!�8-폽�"X	L��V񮩪yqI�8Fih�&|�
6G��t���z�*uO���Qw�� d�xc�#�%�k�^Y��ǝ$�4V@J�����,�	WɑE��>�E�[��d��䯞/�C��7���<C7�8 Ҵ0*�~V��;�X�UZh��̂V��Z Cɬ��D����j�`��H���B�@MwV#��ƹ|W,J�?���Y���$�G[���_��_�U#��i ����U�w�պ���b<�/�@�	k��>���Ǖ0�T0�&y��'	���Xvj���o&�6~�'a��p�[pk%��w6h^�kH�A�$^�̓M�k���U	��4�wi�Q�-��K?}��?���g���Ǩ�� �"���*�[�3�1�K�	�yu��}�-�+(��Υ�B�c�Z�n�>[#�
��)*ȧ����.w��p$����PK1N\�J��9��N�F��u�d��J£P�T�
/�܅��I�!0��
��ȐW53�T-�"��	g9EK�
о����~O�Ý�@�[�5����Q>��'|���s��Ĕ�_n�x�#r��F94ܹ-���]��d��;�&���o��#��3
+!9����tf�4"U�����QD�#�{Mp�tE��ć作� �l����45H
�.���tDꐅ����y�6P0)y�)avS��vw��,x���h�E	Vރ�\!�і��,6i	e�,��Kl�58�r�3�[�NϜ��n"�����*��.��:@�e�^ͳV�<��cEˀ�5�?�@�6G�h�q�>��t���+�ӽ��I��1�cJ�����C?��
V-���*�ղ�A�}R��e�a��?�g�/�.�^��(g�h���{�(�뵷�a��	׍w��EA��p�X�Q�f1�]ێ:%��j �0P#��}g
��p $�����nsbu�χ��b��*%/?���u:t�UK�q�H��:dG�l�*d��������^�.!+�����[#ӑ�����ܣ��p�B: �W��҉5�B
E���Q�'#����ӚWU�u�Ļ����������Մ�03��t��,=�tLؓ�1�D�Rj���SQ�j���l�屓�Ǐ�k@�������=4<w����̋���[r��fA\Qs<��J k���5�u�Q?G�5�Q@`��U����s
 ?��0�iE�ýU�x�f]��ow��*����Ku��'E�:j',��^)�n,_���0p����d��8:-�C)g�7\�q�|\}�*��R~Hf��L�ۜ���X�~��d���e���b�2���P�S��h�¿�Q7q�zBl���e;i��<�I���OM�X2�����հ��VH�,X�&�z�'�y�����-;ުAx�n����O��_�����1{���� ���8F�V�����6��W���l[�De�gz��ed~���U�-�䧲� 
��|3P�bNw�m�Ѓ�ɨ�\�G�ދ���j�rfF���{�(yx�ș�����W�̥ܞ'm�o���ӳb4�_g��&��oh�n�{W���e��t�7OX)�D/ �w�4m���+7�0���ˡE��
s\�k�PT�s��n</`��D�J����������&��[=��;z^�m��{~�����u|Wy���:~}�$7���)V�z�	i��tj��}���m�}&[�	\,KϞ~�p���.�=���#����{1)w�'ޫ�)�yuj�M��YkK��R��i"uceֻ�Զ�Z�n�ɨ�\�>Óo�E��Hst}��i�&�I��C��G��OTJ|t���=��ը��>�i��}�l �>�M�=������H1���t�vawG]�!�w:��4>j,�u�A_���A�4�⫏Fˤ�1x�>:�}�J�`'暑��O�����@����>8���ʳ?t��r����)I�2�?�פ{
e�HXF������A��\�S-���%�|�0�9?�����)�~��lv�	,�y�J��Hf�Z3YQ)���n���I=�#=:.7}tD)��&��3����,bl�E7Ϥ�z�hf�0�8�l�g8��]nX�=N�OU<|����7���/�b�����Fm|wϝ��՝%?�s��h�~U�q�곂���y�R~��\��qZkH��&�)ޛL��^I���pA��(�e~R"�����8���{=��\���5�G�,�D��9.&�����3�)��p��6���]ZuB�o��6���p�Q�ļ�<r�`�"����lާr����UG�Hb������M�g��d`�Ō�(�J�`��j�oA�����l�2ǵ�7�s�l�L����q�����ޤs\��ur"��D�:j�]�`1��C��R�#v
kFz-k��_EOUc�d�گ�]m��֯%�RQ�bߠ˩�������H��������r_Y7�r�u#�T �t �S"R�J)2�k,��J9��/�3hy��ɻ��2-zȤ|�=����ϩX�N���)k����Ǥ�b�=&=]h�ZT[Q�VȄ�r	� ~�]9��}9�ٔu�2������ަ+��`ej�F{���:o�S8[(W���?ˆ��!��6M��0q�%��B �WC'�ߥ$b(u�7t����j���ݭlc��%�x�/�S�K![��ћ+K�L�y�/]~��D5��i>4ݵ�XK��h�����=�ٻڗShӝΡ�U#L����V%L�0N�,�l����拢��j�H҂�K���v�#ڏ��8b�B�0���w�^(��,�e�2�]����]k������l��#��>�3gz�����k���B��e�C[!�~�F�ISѩ��K�w{�Y���~�P�`���=�D~F�+��XlxVHYEB    7d55    1450�Q�ݫ�A�ʧ���D�����R��-&�v2�rV���� �9��z���  >Z���]"ߠ�$�KG��rדN�WC����k��ĚÅ�"�h I�S�,rx%v�گY�L���Ep��u���^��������a�G�r�����
���ļ]X)��[��;�RӈaKTe��0��N���z�x@�G� ��XZ�N��=��k����$T�@zN�Cg��߮Fܯ��Ο��zZ�|�m��*�]Ô5����y�Z�qC&���O�~b��Z�Br�`�14�'��M�|�������
�}��]�\����f�2��Quw�s�kϲ�;��X��Y�z��p/��M�0F��t��u4F=2�E���R!�{�@���ϰ7;�הD�{��S:�@q�MX��[��Ό��/�%Gq59ğ��){[��a�u��#�Y�Z���K�Q��L��3b��<�,\�V��R��2ŵ����I�E?�����6��M�mM��{���C��=���^�&�������u�E'��ad V���~@E}=_��x�o!Y�c��F�RF������(e�%wt���(��/S�d6��:�-���so�Ԙ��h�c��3�P������Ջ .z`���+m�-�vi%����jSV�[CN<��&8��Q�!�5y��L���χ��.}�ϝ��3�h�6e<��Uś�:L�̆�WLӆ{s��!`#�#@�ɢ6���/�ց��lT_GE"%>)t�������rr^�$�5�s/%�������0.��x��l7h��.	��Ǝ���X�=L$�a,�ږ�_��b�m�.�O˶VuߝKlrk{�5A�E�B:C���p�V��1�"H��6��;�@�/x����o䥿#9\�2��N`6l=q@Y��X����߻��t7���Dp�O�h�Ll
�^���tS+ߵuK�`|��,�hwF~�|:J�=b����yH#�k/�9��f�]�S�c�njy_�a��r�+;��U���F��N�$ܙaG�����������W�/w4/�1������Y)�.�\���e���X0��^����4D�`��?ae��1��g����H�P	a���t�[�&@�agFQ�u���� �fhm�+�ڼp�W%;t���}��vzE�^�=8�y�/P&�ʉ7��}5;:�츀ٝn�'�9ލ�cT�`�\��s��]���ҿ;iR]�^�5��n�h�N��nO���b����#�s,8'����]��F�@�Ype�\���+��+����H~�h���O�Y�1�>��SϨ��i)��ܗ�qT����[����}�T%�(3�22AA'���uX�h˵H��`y�O�K��m-e<Pv��q�����Ϸ�u�� ���P��S���F��1�rl��Q5@?�l�+�B�h>T��_GJ��Ikm��/�nd-���	˩����^�3A�߆KU�5��A7�=(��oV�^�����%$L��7V'��q�Ds�`Ei������Ct�ш|�l[f�ƻ������ҤhyJ�v��+�*Oa�
�E�+��MU|�zH�D���Ǩ9��(P�g��]Y�*�� 8�F%[��	� Vj�ĭ^)�@7>fOr�h_�9��t�U�3��;Ήm�N�A�E��Ҳe� 鍭@�/"����\=a��
M�c�MQF�.�F\%��^k΂�'R���sCѵN����86BY?�@���h�t!+RFN"d
�og�,���� ����@9:�M���Z7�x�����\s����P��Zׅ����t���	�a�Z8f[�i���:�:7%�aM,�Ӱ�
jih��{j����;.����\I^�ͪ����* ��[�W��v!,R-63O5�R*���bI.�r�Fe+ 6$cJ�i�A��Eĩ�@c�X�G֚$�?��O�n�~��BּQ��f��|g�`���ъn�+�u-��g�FZ'��B�{��&�Ib��%���֬�(a�
Ŕ|�\��F#��9�y�b2ӫ�I�t�I�Ź��6'{����IE��F�3��x(z�� ��OK6���
6\1x��/lC$�׵?���~
	�V��u+�*b�������9n[�y��-.6M�Z_WBƼzuy�USC������Jѻ�մ� �D�V/�e�dk����]�E�{`8-s�>|^4�k8<*�d(E�.!�U��\�&y�l���	ݠ0�C�>"�V�ɁFqɼ�ő���^+�*L��fFU����al�	݈����2������yEN�U+�Bes���g)65w�t=�6T�<�G��|vu\�����[���CJ牰�TV�~�apb���Ֆ�,�N�{֛�.���~wg��+�'�L��8��.ֲ=�.V�s!���z��K ����j(͡�Z��
C΃p$�����H��ԝf]q>i��Ht��x��3^YJ��g/o� C[σ�5���˼ϗr��e��%.L��M��Dm�H	q�[�&@�S�:¼�ѻG����$���g?M�E���q(��@�"+���K@`�I�۪�:�G��6Vx�E�"R�{�cX�n�h�s]�e�ג�Z�*l��!��D{���b�Z��ؓV�J2{�ۮA�5���z�ʻ�I�v5�����'������v�0�a�7Pvw��.sU�7L��ݪI~F^������Y�b¿��� B�vO�	^�?(�B�s��0���&��1�4n��I5��ok��h˦B�U�n�2p��^�( �p��dA�l�v�3� b� �V2�]�puPBt�ĸ3��7G�T�����͵9��n��B?\��	�RP��m&eA�s�Y'��U&!�,\���9�ǞO��-)c*	�*z�N3�fҵ_-a����CE$y/8���#��q�n��*j�[`�/�hH`�����+�p�,㞦�Nm̷KS���Ǭ_���];s����0��P
yq��8����s|���y�����d_��4!
,��|K�G�|���6��Kd�#�9ׂER���br�хK($QvT� ��O���6l�@U ���HpO�O"�v��}��9dQvrC�&�u\�-qi�\����PF���9~�Rih`;�%Lm�r0�yr�Kp�F>;����އ��d�:�8y��a%"=ٷxm.`�CIXv�Ə�"��$jv~D�sm3�W������4���\�#������g�M�����S¿�JpUv�����=��|�y3��]a��0����d�0���ӷ��8f��1ĝNn����B������T�K�I(gZ}����H����<��t|�\鏫O�<��ގJ���$�p6�CTx��i݂��਀���Y2�NR <��H�M<}�:Kc�/aR��q/-~i�P����P�{�L
���=y��[�FxM_���q�(k��,&�W!��˞��Ͷ��bp>�RB�ז���(͞E���W,¢[KJ28@���y`V�7Y+}��23�(��3���]c�0%X��[
��^F�u�y�6c�݀��r�� ӷZF�M��A��1wV��0[Y�y��x�$Nc�D�L��xr����9e���������e`���
v��Lq������o<�B�~=EwX�T��w�a�<36k#��t���a�E(�^z�#~�8>���` loƕ��� R  �W��S�A��Z����2������������	@�T��a�
����k�lh�Q�Z5�T'l�F���n:�&����5pI̢|~��J�q�{=�m��m|���}�+*|�L����#�ْJ���𢍗r2������+ـi�����s���w,V�r�p2��BחC��2 ���[��(�G�rU,7	4m�Y��T*�����(..��{�Be�^!��"�3�G��@ˡZ��2N�Ҫ[��i�������+��ڋ�(�v��n}*���v:�x.i|xݶ��*Dsb,;�U�ߺ��ନ�f}�o�ϾC�8���p��TFA��+|�� ����P�j6��NO�	��]���h�oɄ�ʍ� �#�ם:e����:q8.�m�T"��@��nCsA�-Cw��\�S��TFi��7.��<���'0v�1�ؽz�kikv�:#���c�3����nF����N�֚e��. ���w���!�v�(��0;�1Y>�:���3ۂg�x��Ӂi�>�*N�z8�fY~��ʌ�ȯ`=�	-����)�R]���#��n^�ˠ�[��50rp{&=AZ	Dv�m��/���ڔ��iC�n�?�Ek� ��k�p��Y*����4��3���7R�+�+u����6� �/l�XY�� �����o����U9�RKQ����Q`)�|	�f&��X�rm�k�"0���y��=K�kR� �d_��i�s��������M�6��C���,��|�	@�����H�=�/�)�d^=e
�A#i�c�t� g)r7ыȒ������v�$=����� ������L�A�@ڴ�s���� w��	�� ��u��xu
�4N��g���(3�\�ܞ�DN2HP�x��*��9� ��)(\/kb9G�\x�eAA_ar�TM�N��#�V/����Oa�#a� ��$[������Z�<%ą����ǐ�xa�$�.����I���bQ�X���9U�U�f}��K6o1��B� �N�v	���nc���������~���)�hjY8(�\[`\fW���ǫm-�M	v��*��me��O3��L���
���ȣ��`����E|�kbwD�new��'+��34b��/�U�UI|�@O.��M�>\ڿh�}u��pOw��s����!�:B�i�?��Έ�{�8&��^���K6�)�S�5�,�� g��A(���V%a�h���fV�-|n��s�P���%E"�a)˛	�ԫS�2�/�kPz;eZ�g��cN�`��~���k9b�C/�R�ߤi�.L-Zؚ`<�>�}pN|SDGg�����x3�˝w��:��0�����[gg��!��D�I�n�﵅M��mq�V���FC�M������._��X���ݓocy���eM�hI+�
�n�D="�*����n���-��U�~Z��М��e�g�ݪS������q�IM�L3�ef�#�N