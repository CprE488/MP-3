XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��U<��*���(�dwSln��t�n�%y�&!��c� >�Tq卖�|�����ɓ�fl���Is�i�Uc2�`j�zU��'�A�0�5tG����|�rͺ��9Q$N�j�
z{��=s(}�,��ֶ���D��uJ�; �ͰlFUk<�𛙢
�p�m�@f�p��h�*�F�V��Z?/��:
j��ˆ��[)T��,� �^$v�q�鮏�{��Z��Ўc�Eg#�ѨgIlAà��dYq븲���o��Z����{��#|�����'qr4K���p�@���k��1�_W{��)�-^0&z1�����H尟R2l�F"+x���z\�H�Cza �jZ:��B���D���S�&a)/�������ɨ׉/񘤚gw]�C`r�1��T�o�z���r=�o.1}
�t�� Q�Z�5�1-��]���i���-U8�$�l�[����b��V��x|�]�ΨFܱ�d��+T�\Қ	r�i�N�S�fR�40B�u�O�����0�q|g�!��Z�;�i#��ܣ�^���(>Эu��e�k5Z��?����!-܀V��q�nV/hr���]BXi�2�ۭ:�J��JbAmG��~�9IbS��Y	�x\�~�<�<��}�h::;�>Z?^�� ���r��J�^��4���1���OR��h���N�b@�iJ`6_ĝ�n�#�L����ɻ	GG���>b\k��uE�9��9�L�����Ao[�qe��фQ3��x1��f�Q�;}Kz��xXlxVHYEB    3da6     fb06y���;C/�?��COfM(Q�����e�qql��^�\�|��3���Aw��w<��RqgFu/`X.b�)݋�#5>��fR�k?���Z�DS/`�Q����@r/�sg��dz�*ٔ�HB�aq�n�FkݛF~wf*���@�r���O���7[S���|Jr⤎j�d=�m������b����C�ω������ ���<\/n�Ѝ*@=�U gQ'7�,3���3�K�\����M��Y�D��t)s8�[�q%�e���GQy�݉��yg}~ᓓ6�1v?�,�X�ᄆ5�e=�<�\h��giA��ϻ��-B����07i^Z��Ee"y6�����frS�؏��o/jC*+���p!��6����^fUˏ?� ����Lc�yL� �: �2����FP�,����Yd��qH�S�Ȱ'��[�����1�^�9��]�%x��U�-}$����B�<�eA@��e���&���p0�r$�2���B�B$阾jS(���Ej���pT�pb��YL��˝�f�p���%GD�[�*H�-�*4
�uT��8Nx9P�!|�K�'���?�$������xXm�3���~�} ��u����^ڹ���Թ�.��A6:���Ǌ]R�:��D1��ґ��΍[��4w�$���BR���U�N�`c���۰��J���E)���)�ds�ߞ,	�$�+?�o��B̗M�Tg�K��������dO{bu�7QP�\44�/���EkϦ��n�m�H�:{>/i����F�
�`�$|I��\U�}���&t|gZ�zŇ|o�G���#k�����p.v�Ď�]�a�v/�y�����@
:���*C��0��|Vbt�>��^��;��[�)Cc���C��/�R'���z/X�8��eO�XG'�j����#;�(�Ԣ�iH���4!)�D[փ����s[-0��%�<9���g�^������b9��ü���1�G�ESD��<Z��5�w�)��2R�1	y��m�3[cvɾ����Ұ�Q����N��;�z�*r��I_��v�p�$�[��1�·���xi��V��\0�:�v_�l6��O����,NQ��p���d�`cf�C{�X�K�2�9���1��}צ�O��"�G���7�QϬF�>%{3 �ӆμ��RK��0R�EJ�Bn����vU1%7�)i�6]�)��DRN��2J*6-In�[���1�t/�U�f��ot)u���ՠ�lV-f�N�oEpL6D��������'_���'9���Ut�Q!����퀍���j�(@"�����NK��b��g�A34h�\�ᖷ�PJ���cB���9X�,��8�p{(�g�)�u���0��a��G˽�w��sC,�z����g�@Ĝ�a��v~��7X����\]�F�˗����v�:5ý���6\�~Y]夃�dՒ�I�@?��F���W~d?zɽX�*$N�|m�5N7c�t���C�Y�ExP�R�좺`Um��Ȩ�s%�w�R@z����9?��rU.�>��FGޞעH*�� L�5!	f�nU�a_��^n����MX���Mr�Dx G�-P�����S��q�
�1c�ğ@���cf�1�L�D\��h����r �x>��;���e����M?4�/^-�x'ɩp/��'��&�܎MByTi�M������O,����W1��#y餕�_�8��GK�R��I?E�UY� #V�����T��qiˊ�Ņ��lSҘD;�U!�����u,2~��� ����~����i�9	b"ິ5$:�]d
�����dz�s�U�;$tZ`b���h�H�����`Qb鴖-|�N�'pu��5��~����%b��zCǱ�ʭq�	*�~E�����\�b8�q�Ǡ�0]ېMj�K�R���2�P�s�O�G"�Z�� �k�( _�M��ե�v�s�/��k��|�qmu�i��#��&Z��H�+��<̆Ⱥ����xk�;�嫼�k}U�*����W����Ơ�
|Y�5z6:m0��ϐ��r�5�$�R��#��`���R���Ӄ��跽��ش%NVG2����˅IO�p͖S �L��T�I7o�@���a���^2��i5��)!�?97���l�G���a��dp��/��L��[`�Wl[�p��'ĪM��\�>�e������Q�+��ru��bt�d.�˒�jb�(u/1��/YN�.��$ܥ�4��<�2j��i���b���ץku�SQ�!a�}&a��P(��T��1e���F禄�AX�����q�2VfP��������ثdJ�kRPGc����l�f� ��>+>dX>���+��&�^/�=��G�ӡ$�Y�`����mWӺk�4pr�ZL��죗�$Eoj�*�*��}��,B�N�k�̑�� �T�_�sez����6zo$�y��/��ah�I��ۺB�
�G�l\�-��L��#w��A�KF���C�}��*Ħ�Tb��,)��J!e�4�xN��A�e��`��,���nL[�����Ѽ �GL��і�H3F�0�J,~���`+Z0F޶z�\#]�Vi�6��S�X�e/��ZVw�l)�Or=Y�#��Ο��P�.?����9QSğ	v5���W����*A�#����4*`Ii��	έ�/��,2�7,�.T��T���q��f��T��.��T9��H���9���:�0e���cM�}���hU�s=���v~�ЄS�h�NZ:��"� ����݁ݮ����o� w��X*�{6���5I:��,���/%rC�4����_��(7Z����<�u=pG�nZ���o���ؓ�X�=Ŗ��z���Y�O����N�!�
�
R��Y��<������5�1���|�6!�|���ܘ.D|�0ݼ�kJT`�=���
+]}e�������S�"uy��(���R���M��67��}S��ߜ<��לl*�%��|����Ҭ@m�����.�
�FUR9���z���U��LKi����ۤ͡�ѡ<Z��39B�]���Q&o�sBLe��)D��Q�L�����\(�=N��|K�-��- LFVh��O1!�*(x#�{Fj7��DS;p!��4���"0�cs���b$�H�O�Ey�����f�w�dv�;��;��7� �3e<#���a��yM�?-nD%��d��",`�}�|5ڄ�Q)�d�[�T�( �+P8�sIp*�M��5��5�8�U߄'��J�S7.A<ǧU�	QO]T���rM�1�Q.˞�d�g)W�Ɛ+AV��.B3<Abu�]�ay�s$���̦�i�s��}a�)T�H�O��Z�'A���6d#~�y�1j�~rQ��
5�}yM龱Y9�/'	r^���c4�?S��:9(׭�zW�/2�����������CحmBɣ�,6c�b�(˄t+
��� a+s����a�P��,��2.+�ŋ1 �+�>."���N�D�;���a��tH�k�ž��
$1p���N��[��Jb�B4Y 1������5�,��g:����fV�	J��x�I�s�/+�-R�V��UHlt߀)?���r�W����)���O�	c���b�orC}4�9�ôW������d�*(���(}�$�������� ~- r���L+���oz��r �)���;�\��ޓ�CN��z�4�P~	���4"}�N�V��N�y1�m��y0���F{#��w�"7p~b��tK��A�:AU"T? �6�Uם}���E���Ϗ���h5��?���"K,��r��;�Ts9�F)0�}���y���H�����L�x9ba���dM���
��f���QH����
����T=t�Zd�����5)N���0؆q��1�|Р��v|���