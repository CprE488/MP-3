XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���VVGyzoG�Zh��(�_���[�g�BJ{�3�Y/�o����S��@ �r9�HQA=+9-�=�� �%pJi=�dƔ)��`IUrOG�v'��9���k�N��V��!�=�I)���l�ᛥX|��ތl4�T5��m�g����l���H���7��$xn���'���I�c�%ݘ���qB�����Ӑ��i�^��Ϟ�t��0ѫ�5[�O���J�;��8(�Dמ�%
���20�`ЊH4��2�*���gB�U$޹m�����Laa��l�]�B��:|�N�e->N���_#0�Zq�d����`؆#m��x49���B\�'SE�,�SXG�O!��4i�����o��[��RD[ƪ-�� J��y�}���[u^�[�a)���k &U��akL�F�pfJ�O�d�T:��h�:u6_�
�bѼ�U�MW��q��B�Xѭ���m�w����� ;y�ʲ�1�7����2|���=��}[�kqTx��E3`;�j���ᓾU.<{G��"z��
J��@�-���[�)��k��)g�m��s�<��B�"{L!2'�8��	2%։0{#�� ��c�GJ���F(m4� �׻ʺ��[9�]E���ӛ������9���YAwDm�#�L%>�����񶤲�յ��/\'�qz��W�z�r\s���"e�UFr�B���!6���.@NbIU���~��ҕ�S�Y��ӛLux�1�^��!8{�*��ᐯ2�[��p�����o��٬69�Ɍ�`9XlxVHYEB    893b    1e30���.�vੁA�Ќ{���{1����H�Ԋ)�{E���pm	�����)����1J�][��pAi�����hW��|D'����[Lֻ��"���*��e�!��9]�� ��v}z,�Y��{]3�֒<�{�uOT�Au��>��٣ⱟ��>~�}�[RC�Q�_�����
�P�t��a@��u[����8�h9Ո��s�� ��F�NMG�O��hIVʟ�V�\��BlL\ӹdvG�YI}����+��J1�h� ��\@��C���"V_e������$�J/(���ܲ��̫ܜ�_�#�2RP���h�q�奟�Y���iO��9ww�+ri ��Rڇ�sr�Bs,�hK��<�}D������fj���-LjШ򼝸�*�]���0h4��+�Tm���	�_3���UN�o8�
����h��������Xeu�Q[{ز>b�����q`(�ji���;�Y�@�!:Wb��;�O�D6K(X�g%�J"40n]�����λJ� -)�s��XP��{��A�'��M�h
Ȕh�L_���"�H��?+S��*U/�d�࿗to��X�Lf\�g�kE}8owt�ۄ+n���Z����H���0��A�Y��r����|��l���'TR0eB���ϖ����Y鄒x@2&:PI	W���%f*TpD�J�E��.O��bpe��������l�V>T������ДN&51Nht?%_��B��jPy��M���CH�m	�ү��@�[�,�� ����r����aЬ/oo6�e�>�y���4E�n�1R�b�q`F΃MJC��pb�S�{[_Uc�������<�^q��rd��`�Ci�>����@1	���g�|�T��J�q���	�G�.�;>��������U�~ϖ�._��N6�_�)=S�sM[��.IO�*ޤY�LXw5t��~�d�`iD�w��XR��.Z�1f�lJ��5!-�&�%-~�������>�{DS�� v1���-�Z@p�|�aZ�ń#�cA�gƐc3R��o��q/��H���9�Y�^��^w�6��ސ݃��9�Bc�h>t�T�L3zgx�`�<�V�VN���8�Jq��]�]VvN�ϷA�$���-�zw���g�	�]F�Qt�
в�w�X��5���h[L��S�贘+'��6>(t[�2���f�n��5p��-��1ToLH!�m˒�ưZ�LJ�c�]8��~�x����.~b�5E�[�A2|瀔2��1���#�ިbC2#_�N/+�2Gԣ;.����ݭ�?]�zmY�Rz�cQ13���_��`I�-�t�����:*���ψ��p[ \5Қ��d&)���<̐�7QE�7�#���!,P[P5���T��>�p"�c�:�aK�G;裵�H\8�� _��3L�.����>)�B�mL��K����ϰ3T�-�<������0+E��DF�vށ�F�+ý5��3�i�مI�"r��m�Up�ҧ�
�Be�HB�k���������B3���_c�?�Dm�.7�����1�d�HŭY�^*�*����\�C�
��M�3H�א�Wߦڤ�@��&����h�]b��Gh��;}}�0���q�-�;p��p7�&�zAȰ�8�y`�B P$��w�s<���i�\���u�c�.Z%�M)�a�4����S�4+�{a��0Dv�K��,�,�I����S�����3E�В.��H!4N�6	.ljp��N&�X5�9�-n�H(�^j��C�L�*��^�3����-8���K�gUKj�)v9��o������{)� I�lՇ��ݺ�&�ї�[�沊��B�Z�O��H�hhg.B�O��Ş��@8������u<~]hk��Rt�ȱ��՘}��U���Q�3���nk��.�S�X���&ǜ��au?��3�m�r�$ ؐ��pj�VR>�3��5 ��C�+�u��Qd�6O�r��l-+lܝ0���z�=Ev���c>�A�z)�_���	�J:�'������y��EZ[q�EGt�F޽&�B2���U�;���f0�M���d�Ba19��o��^����2�:����{�z�p�AW"Ie�[v��YLd�<.���	\E`���	':��@a{���X��u4����)� �0c�����>�!�<�'�G�#��H/
���[�Z׶H,G �%�t6^���ך�~C=C9P�Z�,�Be��-����*ژnF:Uvݽ����gI���c������|�=�uP�;��9Z��&�FY�,VC�_\�����u�y� �^T͎Ѱ�;�t�r�i�-���KՌ�����#�߫w8�X="�u[�K���#��9�>H'3�'���������a�F�c�����_�뤰y��uk0�t�9�Ӈ	���n:i6�M�T�B���(NǨ��H�MѿHv;o$%�W�8���Ƿ�"�9���,[��me��]洸T(�y��܀q,�K�m�b�E����?:|C�ĩ��WYL$ݰ#lN=�T�����zM�5i��j��_C5�2hZT�Ұ#V�ٞkf�/�X�*�@�C�pT	L~QׄX�\�|W�~z��/�<�F�	.���+����5N,P��aУ������Q�D͘u�L�}!$����K[�G��f)bɊ���Y<Z��2�H��_?];h��e��[�P��}Z��0sR�l����r7�.&�le�3��6�ُ,ф[Vg׶jP>����̩���ۮ\����E���֕�2�i�U�s��X�KV�a3��C [�뷝z��$����U~&n^1Ȝg�')��;7GDenu�q�FlҦ�U�K��i�q�t�Q��A}�y�-��:�ߴߜK&ꅰ�4)}:�*XBx ����=�=���oJ��cK5��'SK���xn���Ǚ������i'�7�|�B�bju��W���:��|hg�v,O���W���\�,_K�2��&F�$�Rz�ڒ���h�eU���$��3���̞�y4�c���$��3����J\-��5J�L�˔L b�ʻ@j0֐�.���6����K'7��:?��2��"���JŃë�-��ƼN�"�]�55�痫C��"�ȇ���<l}�Z@1����4�H�\|��#IӠz�⭇w>	/��A����#9x�̂��wX�V�i��_9v=���v�?�"�Q���i������I��Wd�Mi����S���Hc0���c#��Px���rJc E�	��,T�m�6:���!����L\/��e�T"��n�MP@mA�w\��H��ۣ�������y�ezx������֓
[Ý��E�=�����+���/��L�:��0�ڍWԇK�J=⋫�jO��TB��6��Y5�=F�>���{�Jf������Ҋ�)�L#t'I&���I&ߊf6�a��<W ��س�o6{=Sֽ�"V���a�O3���)Y��H��ӱ�Q����l��b}�lx︞�f��N.Q�i��KH��N�0y���F۫C�j�5�n*�𹾠l��	��	�(���VrZ�"��Ȝ.���7��}�AG�Q�8C��<�b��
 	n�a��������o�w����%KX���A�&4�6J�]�w����/���a��o�~�����N�zqc�w**�A�O��x�yU���;�R/e��ιI����� 7�:k�\!{Z
���i}Uh�J���p����+��$��[��?�T�cS���,���4������x~�5�Z=�B6hXv�����S(�q��zt����H<�w��߅���K�>[,��U
�S�O{Qc�U���ڐ�x>�-\!]\_�zW
�:GD���0P]f6�)![��%n�פ9z�U�ءU���!KI�`s:���n���i�W)|���Y�s���!��OE��B�@T�S�y#�r��W��^���8���N���X�:_���A��{�ҝ���^�<��x�t�A�vJB��+{n��o�&L.�"�(]/`^�S�+��2uI�X
�Q���$���.�dj(L��bbx�	�Xv
'��B�B�?}8$ݶ*��>i���C�āIf�5=��zj���"�AvxJdVl���y3��Se?H�J��cR��� \��g�/n�x�=�e�4�U˥"-��C�Q��R�<+B���j��*W�/L9�J��V���!��'�I�_�n�,�{t����on��P�&�&�=D��P�J��S�)h뒽���r �E�����߼�u�1�<7���h<!�G�����qA[�Ə���[Zq���b\���+�I�~'ˡR���g����c8�Аg%\�u��
y�8����!J��P��8��pb~���9r��繑��i�)��Ĳ�������(�z�h�X7G�G�ֻX�8�"�Zh�-����3f�3��$�F�t�������-.��� �h��Ļ��@�7�u�Q��:��#�m��*	��mI��!��:̸g��C�ذ�%ܹ��6IU@NEQ����!*u8� �c����S�1�Ɖ��k����;��5ʾ&x��@�юH���Y(#��oZ�y�Ɩ��b��1���X/�������ݾ�%B�z!�
҃w�ZU��l�6�g�w �?�:u7L����_w�PM���.�E���Z�������|V�fA����[�.���s7�xy�ǌ��&���F>����*�'��a��b�ߨ�~�e�'�-1�&Nt�|�G&���~�<�8���<Ԅ�ߙ��w�;�d����hA�(��׺GTJ�Y� �򣺵��(�*y�4��.1����B^*ԘFȭ�m �_H�v��ޫ���\�������F�*��D!V�gs=�Zh��.�
Yu�@9�J mK�71�5�a�^�d��%���њJG9"��J�u2*J�9���J	f�X0�7LӤX�<���s_�+WWƌ�� �3%����cvNr��.��n�^�jJ��Wj���2��S6�q}ul�2�u���G��0����``��j^Mq,_���3��o  (�P;F�kRf����p*X�������V�
�n|�f��u>R��DP�ɲZ���@�4�0���||�P��h�J�z��Į,�݈\T�]�:	��|{ .VΣ���=�W��C��p��$�S�p�.�h�~P:�VF��u|�Ӡ���HA���ƴ�U�()�+p��2���ǽu���8�!�b���j��y�[`@å�S��jU>Y���.q�S��27:^���Cb��t"�� ~Ƅ��(I��J� �[u��:���o���-����&��Q2��sR���[;FC�4k�����r�f�S�ϯ�Ùр/�=�Hu��p�'+���i���1F\���D�����gQ�x�}?�Yt��G�^�7H��E]A3Z��!
��������2��S���l���bX�%�~����h�ˤ�q�zЌ-���{MQ��mO�`����a�mb�/vR�J�&��^ԥzQ���0Jp�W�Z#ğ�����>}S�KE߲�Ǖ������51�ɞ�N��:[څ����5Af���ZL���o�C��?���}�RתO\�3i��LA����T��"�ig2@T�'	���s#��Z�X�	��<"�L��c�]ͽϜ�����<��=V?Uvj��ϵ$7��Q��]c0��s�ƍ/���m��5r�p��c_df��)ɯ�X5����%L,WFK����wu�Xl砥o*����^���;�k^��D`���R8���̰���U��ycs(Q@!���gق[�7�����dg�����w�Y�
�O�-e�9p��Ԙ�.�]c6Y���ܣM���e��e��N����A�J{h���*�*-�m��|��-th��a=z[[)�d��"�/ �KUM{��R9��Rl��q�.�{�m�NedB�U��鮹�!�j�U،إ�}@ǁ���PY ]�>H]\}�[�zS�ӥ���H �J�vw�+#�*���Ȼ�w"��#��1@9`͜�����c�]��K�t��K�`�Q��n��d��D�B\�����2C��F�x%��[�H���9j>�h9R���rjQ�T��$�)
M-~��7��#��ښ��1
���DL2x�

�y�0q�>f+Zd�c�5Rq��h�ZS�%��D��\W�
�
��/)k	]vNu�!z{�Ƞb�t�e<��
�$vf�A�0�Ri�{�,����W��(���X����F���Y�˰�����s�/�m������+��e;Y��;�r;��&)�B,7˞S<�Vf�F�l>�a� ]�����i)��􎌁=w�m�l��s���NC�+��X���%KUI$9�D�߷ɁկSO0�p��?���tD���?f�^Y�ݛ����\4��%�q`W�}����j=�G�7����1�p��*�&Z�'�d��o�C��<\�!��p��gWO�W36������In��~�$��/!��A�j�
�ax�YnYK�A��i��q���qk����`����#�m��lJ�^a2c��U�${�%Y�0hj85 _���]����^ƍؔ�_	ʪ�3.�W+ll�U���8].��+Э���0U<d=������
-�|P��9i`}��ҩ��7WHuL��������:J�W.��ǡ-�O!(x������ȇO�l��p��5���@��c����+s�]`�x���A�L~@�9�%�4I)�i�ܩ�o�B�uʧ��g���6�����������2�$�jC��R��٥�<��$�(��+U�~L�����Dб)F�$��yh0�O�V�d�ڒ��j��+��7pv�n���1�BS$���~���F(D��,_�t�)D��� �.9V7���b�<CSJ9�z��)B���9Z�@u�B�ˬ(,��Al�ӭ�XI�?�b^&��Yy>���s�vM:��0����`�su���-獠���U^�՛�J؞�� ��ꭲe��^���Q9¦�[�9���@�W׆*����9H�N����c��O�,>#��I�B��x<�*��F���eW�w�Q�5�zi��^&p�m��N����j\�� J�U�^f:�$��f��\�%�o��Q�|��9<-3�~��%|QG��}�4 7�3g�1��8Ɔ3��1�+��r֕Ⴡl_U�� )2e�i�:����(�	^Zw����4J�L���(�#��,�r=��6�Z_����}QH��s6Tn����b�XYU
J�ua�(_��v\t�Ѐ�@u�N�ANU�b�LO�&{f�7HD�h��%�Q�H�Xܦ����j����T�ֈg��Ou=�����dLJ$۾��d"�K�bZ��0�Y)�kp��������1�#���-ʘ&��􎜽�������_�d�S;���bK^%�d7�K�x��	�����5FC_�rA�,;�	4sN����7"<i�u��H%��備B�0ٯ0�,�M��\�E�宂~#]O,�_,��{W�� ��@�8�W=��cc�Ƥ�ڊaX. yi��ѠD�m�h;����Q\f�[��ۆ����B����[Pc+�����6rV�@��"�Y�po����"B����܈Q~ѫ��"�Mz#��	�}����Uk����>+��c_Wng