XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����3����@(�v��k�U����{��	z�C&��S�A�Kb3�2D�m�WԎ��ڛ�g�ә��[���z��N���8�����&|���"��D7�ް~>*�g�SH��6|�+n�W\)�4��DNp,c V���A���<�)��M74�iе��!xt�vw :���y��'��K�I%������o���t����a1`G~����ٙQ@��~��i�f*���ǽ�7�B@�IL��l��'|h~�>����׍�M��8���|د�A޻�4VjJ1��#
�^�x�TQX��U3��?>~��a����i��zE��^����PA�'����;���9(8`:�'G�lU]�޼�7�W:/���|K�ܳFm�ƺc����*d3��3a8N���'l�1�L^A�\�����Td��ab�3j�m(0`'��]n�xz]�J_I�r6WtD�ޗ�����O�S�Ȃx�̫�,iv]�З����M��D��0�@"��p�$9��ê���/!�L�,�1?�f���O~R�zG$;��P�ii��h��L��W�T|�ӺuG����o��-Ro����ٚH[�^�wG����OE �b��Q�dD_]��e�N��2$�y��8��\��J���ʶٗ�.���1i%�i���ZW�V�&�aW���<�����������<�T��`�0��rm���Q��n����W;�ћ�8@���7m�p2�c�h+�*��Q�F|�XlxVHYEB    1a34     990�S��'|����CR��aKH2�h��qv�Y1U��~����[��
е�Rt=�;�d�S�+���b���z�e��C]�܍y Ӟ�0�stSF�h,r}q���;O�����g6ɠ�J~)��2~^{�Mg��/<5FU��Ц�a:����m^7��W�����T�$-��ܞ��;���F [���Ԃŧ�z�${c�dYj�x�	cpv��ѭ��v�<�����Zi�Zp�b�D���}�����ĳ��vït|�����.��l�R-��H�&����I�G/�*P0=���r~�#����5ӟ�ӑf;��W,�:�u�)����D��-�}�ⅿ�y13�%-�-j0'��`f_�}s=�4Gr(�S`u����mVa�c/�S���pG��$,�RK�����V�p:�'X��=8}��B<�G�&^��[�r���Ҍ"F�(�Kt�<A}Pyʯ�.������<�;�#�ɗ��c�������\��H֍�J� �\��mL�G���،�>I=�"�����'q���<����u����qI�](���y���c9�ĸ��2�G 7���y�3}����pQ�A�Վ�I�FM��bgC�+K��%��ts��^2	�A7]�l��=`Ε!�Pj�J@]���6Sx�じ��[,B���t0A
hh7��~���W���zg��i�JXt�.���x+|?z~����,���;}�������!�q!����(:�՛=�d�~Ա���d0�)�n�C��H^z09c�X�߫����,������]/��#3~����I�iLK��N$8$$s\��o}9B��[A$��xޯ�@s/�@0Sc��^q����7����$2F[+�O���Xp���-�`���n��M��]��R�p�=ިe�"^���K�V�����tG����Y����=����iי|�W��q�C����|��r�݇Z����(��(E�H8��g,P3F���pI��xzo���<�p�q��I�!��"�NZ�Bv��QrG� V�Ʌ93�Y�Vp�h�(Fj�ѿ����.AWi��:���Kɥ���2����e��ꫠI����
� >�/3հDG�� �ͭ�}�úP�K���C�� j}{��I���52�ʰ)���GZ{���+4Ha�`#�U(L�h�Ai��\.%I�}k��E7QΆkc�����T=���?sǫ�Z�RX�M���(��筌:�n(GA�5�˹�HZ�ap-w&�����3_8ɠOK7�w����Qn���p��0��R� �]�������e��٢ٻis[�\'!�:��6�x�R�e���W[~y����l��]#��u��,��󞷰��$�����"/.^{��{7���*�s���J{����������d)�)��'��4�u��Љ��~~��<�ݯ$,��Ⱦ:�����-^����C��z61џp1�!�^#�T�Ƈ����c��R�.�����Z�R6l�0H�--�$� ���`����c�f16[&�&�H�0�K'�du85]�R<n��hH�3x��y	v�=������!��g;ozI|�-�Aڦ�4�"#Mp�Y��/o�+�w_7�nl֌�P1�$�(���_�"���'k���>����2D#U�uJ˘��ZC�Ƙ7�/�4��Wz��I�p�k1���s�o�gu��@#FqVγ	��_O���{�v��S�6$!2�򣧘�O�@i�'G:#�(�+_p�X�������vʪ~I���'������.f���lc�2u0ǚ�G8s�����\�9�0�M���
����f��i�_�Xn(V�7/�����w|�؀S���(C�$�]Ea�GԔ���!Q#[S���k�~Se��ni�	T�a�bu�5�b�X�lX�t���7a��,'Nt-'�b�|���; �|qN�[ Tn��,�*�]�Z���gy�� �+������,�R+� �l]�6h�k�V��v.��i���_[|!�/��/���y�R>���C�8A����LHGT�%�ToŸ�e������l;��Z�-N�˶dܬ�\F��",��#C���/�S�������`U�3�@tfҿ��tdB��i"�ۼ���� �	*��~�TГ^|tO�Ycg��.7{Ա���F����ɗ�1��~2��v���:��.�Z�;�,ָe�5��cٽ��I�	y���nK�?n[
t���a� ��	1/	�X=�&/_�-��蜹ω�2��G].�jO-첈��]�$'
"���j3�bgG��X�^��q�����!���0����_�$?lj���]}�g;+��d �AƁ����&O�eK�n=�K ;drvy淼B�1�2�vE.����V%��� �7w��$���M�'���