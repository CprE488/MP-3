XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����<�����2�~�e���t�E��O6FdZx�]#��|����̯]�G8s�#{���~���yL���H��>x��`T�z;`�Aܾ9��A���+9�w��	�1�A�g���J� ̇I�����-��n;�2�<*�Z��c�p�ϣ �*�Ǧ�cB��us�qJ���{g!�!��2����ˢ�����9F��&>6�$F/���x���������!�SXB�Yr������+�~�o1�tfT�8 y�ӡ�".DD����Q"�T����Nx }��TQl5:��.�S��>Ogc�#�r�k���Y+�ov�P�seXh���jeг����RHȡ6b���K"�#3�o
������pI��3������豐�äڭyf0���??bI7��ƴ��a�!��Y��Ǣ_$����mm��;����q�cd#Sl����"%�~�_T�ORw*Y�wV����j
J�;H�/M��8��k�f�Hꖵ/�Y�H���1v�c�e�/q���řo{_[��.��	;5+�?�I�'W`��.{@d��-�s_F�_ǫcd��"v�р_��Z�ª1H���.�ߗ�ˬ<7'��:�����Q�xL���=��;�� �G��z�82h����i�����^ʺw�
�Y|l�s�� 1��6�{4�
�g8�����l� ��y��Wi,M�i8Y�;��	z�9V�!�����k9v�W��𵌅��1�/�W|6P��K'f�6e�t&���|K�Kk�w�@�h���XlxVHYEB    5d29    1390��0�s��ȃu;��\o:H>����Ὑ�[���,\�QP�e2�t?c��rA�>z�&'����^�2�)����r<A�*�%�B���I�
+aO�������b��&�3B��J�b��g
x/J�����]u��<	[e�c�둼���ؓS��1�~�������~�ơ�hw��"�����f��-��D�6tXU�u���R���!���'��K��k;��W��8�+�͹�WQ��bx:#�%��g����n���f[��Cq;���4Y�Pz�r��dhZp��!�Y����E%��)��p��z�z�_��1��������rf���(���A��K�������6Q�������x����!�=����F����Ķ���*�{ֳ�#f�#҂��8;�zE<?Uh����E+�1���{��ޒ�ݬ��u���Q�z��8�P��[�9fZ��QML�zW��Y�EG��߅�7봗31]vm�u f:P�H2%W����qM�N�L���%쑿�N*��T]~;'?
�R	�C���R"(�7��{�	���}��mO�^<.�5g*U ��o�+�{�k�z�=�-RT���3��cA��� �q�\�~��t���� V:�-� �օ(w~`o��6�	� t�:,@+
RV�|ˌ�&�ñ�|�p�u�{��ZQt�B���N�������i?�q	�y�S�W}M7�ʷg�R��Q��Q̕�'�	7�^����j��_Z\����Dɉ	�-Hd��Ų A���Ap���$/[�C����H��C��U����!�C�s��9{9��@�	�g���U��inޒLr�CT(P�#[�nm$�R4sL"w�>��J��"���HƠb��_d�����L�[6��#�K����Q2 �I{�t׽���D*`�t����xJ�]�~G��׌�O��g��R'��	n_�$I�f@S?��ƀ"6��)��9�C���^\�������U�\h�D��U�8:`����lB��j�w���qM2�)> #��.��#� ���b���=�(�DCD	�m+b1��K���Y��|��bq�@^_�ü^�.����~���y"ZZ�IG�t5�����>��#Rnz����:V��ѽ�2*j����D<V�)Q�m��p�޺�%�����m5�f͗�c,L��	b}��"�� � ��a�3�ݴ�Ѫ2:��_��Z��H����=*�U!�C�A�-�`qmyv�5�HK�����ѻ.�3_Z�rFۥ�tE���{�2��66��-��#7厼�B�H���]��md�~OӀfp�3��|μ�ܦ��".�/L.|l�ަ���T�������_t�t���g��0�?>��L�q�4�\5��a<�PENQ�gd�^x�yDX)J�ͮ0��O(��ho|�Vg��7$�Q
�\m�����P��E�;�`C�E�MЯ�罌���߾�H��p�7Mv���
��^^&�&�ߔ�>��@C�/#�;�8򞼱�q;�l�M�I\����}v�]���Qa��4N&)����ۅ>N�0A����uT�>��=��ƝY�$�Eǲ�B��$+���[8W<�It��JS�>��M�c�Ю���!D5���3m�=�ye��@h��(Ȋ@ߜN���ϖ\3�\��\����A��������o�}qc����³W����F�����W�EN�^S�xq�C4Àڴ�Ԡ���fnx�����B����/NM�m;bS����&�ֺZRU'	�y/b��O�C�ٺ�ϕ��.NđI\B�5gvg�C�hS�{�`��7�5�[Ce
��鋞��$d.�mކ<E��9S���@DV�L8,��eÐ�~u%*�D�h�d궕�=�[i�P��|��dI��6��t:��\�&�ȪN��J����163j?QA��}�̢.��@��mǇ�'~��҄c��
by�g��=��T,H#�e[Ex����X�A����p�ʁP��^B��Ӎr+��	Qb'�&Y��`�Ѿ�X��������3����c̠��]~�I�-#�<<@K:}N]��8����jɛY��vb\~~�T�����$�A�3- ouiZ��#����̯�)���i7��t6�E�;j�0�Lŵ~7#.�Yb���E�=U�h_i���P[I�PJ��,��(2�����p*%���x�ekF�wj&��Ģ���r,�Cx��ؚ���8/h_���̎��UmjxE����s�S�Daĭ����5�V��7�v<_dCKU)L9U�z�\,Ota�(�$�J�͘��O?�# ��P�jwud���Z�7�w�! X_�T"FЮ��ݝ���T�#B�b�pL,$���8�G[q�Cz�S�y<u	z3M{�P�X<CS���V�ߗ��BЄ}{F�]�X+G!���2#�
Z"�������6�K��3���T)�>j|u{�+�^�L��R�j�2��|�NyŇG�18�]~��b�$�e�:���_����$S���H���z�䐤'ri�VSj�q1�=/��_�ߠE���n4���V�\��bt�r����a8A�~C����n�B��p���	r����Q{�G:�P�,P rA�����o�c�H":�*����FĻn��^o"����� �?��ÙP�*y%���5�g 
����e)X򢰜D�#��^��3��De�@��8�K�&���ӭ,p�a�j��]�7i*�NP�<h�(y��LG?k\���&�*�����E-ޞI�g�#�����k@t�OSv���\�r�+]�ȸ�����xk��O0�=J8� r6�<o�o@�9@[���Ω���{���<��v�D���x��f��;��ғ���Hk���f�#v��G�Bsp���j^�)��WnWQ��ۮj�ٸÝig�-T.�����CF�{�er,�������N�W����\\���s���w\l֠��AK6�iߡ+%�`U�2�V�)xh�ϏE�~�~����.�|�[N/��V߷đV,�Gi�hH��N+Z���i�K� 	� 戀
 Yǻ�>z��U;�u�J�&��ԣ�����!XSE�40�nu��Z��κ�����u��Wʷ�U.�%%/h�v5�����՘v�Jk���X5�֊,�BJd�`,����=/o��/p���`,g��-��I�f�:�#<0��Χ<��j�`�cz�fs�~[�?�����b`?lm�/.w8N��<�16�����7:�6����O�C��C;��X\k��Tіad|,��R��/�g5�X����o1	��I�k/��M�t^�xEbr��/T��.�೭yB�B��Lk[/%�C���o(����S/rG:h�X���Xٯ_��
�f�横^�at�)#�JŌҕ�1��o�
-g㍗�{�����H\����2��ܗ�GөoW*8Uђ;3���3��X��w��2�/ /Y�	����qBT�V��&�
#4U��M+b��AD�����F�"m�{�^X�@)�.�1�Kr�ٍ�����E^
��bѝU�҇�S�K������Ȅ��%R�_痪u��� �>�_ѳ����J������8�ix�H[���o�U�ꯂ{��Y� ���א'@���Ժh"�G�d��[GG��'����O/w7�f��{Z����4�����l�4a�-�4�᧱6������ ������?�ܫ�ٙ]�&�L[���?����+;���Ck�������Ծ�6{�@�҄�T�Õ��NŇ��Q�ܠT3z�Ǆ�d���ƣrR.2�,���u�0t�4������V���2��t���,���bQ�%6 �&�ٗ��Y9-�;b���H��D��Unc�,ͥ����#{�>�?���}��}u�����F/�6&2z�)7R�����n
l�D�I��*�f
���(����h�
��/+���z$&�e��������x0Y(�3e�@�o�L�kיa����gԴd�9ȸ�|�9q��(����\J|�s��f�~���<n���E0�b�ڽrm���IMƞ�^$�<$�2��a1k.��H���w}����:�����6��-��ϮU������;�C� 5��#�|c)����W$A�M���̊׸���,�﫴9vu���ĳ�|E�̓�,�Rn��qK�R����P]�4�+��~]�s�� ^0�V��b��e��$�D��=�W�7A�, G[ʖv3��N�~Lq���ے�~̬�D�&��>x&�+V�&��h���	��w?��Y��b���	_nEm�Vz�#8��v"�w�`3ƍ� ��^�z��a���J%�f����H5���0ʵo��CF~O�h>Lr���ɱ����C���L�w��<]-��C�^���J}U��J��,��nl��?s����������۠�a�~�T�`�![D�o�z~�DƳ7.n<w[l0\�ɕ�Z��9'�ܿ�g&G�$K�m��+����VfB�p얛�)���jr,)�M7�������� ?�u�n����ܮq.�~��!�w0��	��,�ۏ��H��E�0�E���9=���iz��ufAY�/'|=�5:N ̳��Ope3i�pA�z�I2J$���R���Q�DYlyW�{Rղ57;�䊖�V�jQb���9�Т��f�&���t�:����������ӵ�G#B��irȶ'o5�<��`{�0O>*Z�P�	���h��n����h2<-O�YR���D�ӳ�(*g��<�MM�o\�� �s�Ws��*��)%Xh�8����s f9"� ��o�h����Da!�ⶳh�Pd�4�@3�S�>�ƐYb����{z��$��uW����(�L�{��'��Z'�G6���cph��siYMu-5V�){/