XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���N$�2��;���!GC�R����k�-�M		Ql�Q�Cq��=�Ц�-��"����?O�\�D�
���s�xuK��+���E�y*s��@5W!o�]!Q2�����ິZ!� S�p��< .ڇ��`�{��_�ݏ���^��`�+
��~D�$]é۶��|�fy-��W���-���#^�{��%���No53�9$�X���- ����\K�N�uv�c]���)�����SCK��3iY�	t1�L�>p$0�v��9ΕD�O��L�|�����W�D����/ �Ǡ�PԵ�%��!��(��n� ��x>p���x��"ع��EI?�'����+|�wF�Q����¿tIv	':��/E��ч�)��6l���ȔC4:���8��k��
���9�a�wE�X��O�~���!�
��i4���R�w�V��6���܂Z�/5� X|c����L����m�]O����m���F�������p�}�'��4Mh���p{���D*�h�w����O�v�
�]ճ�%���#�~<�s%�Z9�ʔ��b���pdU����Cv��״�q�X�چ�kpO������Ŕ���f`d��*�6�ߕr��}�:s����8D�"G�(�y"(5���9Ϳ�����\e(��#Ng�%$9w:&9�����8���:���ٺT�*�0��� � L�PK���ϡ�U���e��-By�.�!�;g�]�_߆�e\A[����X,߈�"�Z�'!��XlxVHYEB    fa00    2040�tI�W�vŇ��f�����'�5Qh@F�a��m8��^�'��d���7	��������$��a=�'���1������,u���zI�.�uv��P+t�P��3�ț���l�l�&S%�@A��h�v;�־��[�5����'�"Ϟǋ����� �Z�8�u�$����L���y�η�`?�=Fz�m��u"�'4��E�I��|G\i��?�h�"��W�Qw�(�Hp!��ز����da�0�K,�~\Y2��Uz���`!_ͤm�=��[C�Õ�,�G��R�}��u���ıO�2'�AH�*�{g�'���U��ۑ����R$�TC��E<�<����i t��t�؟(�:�O.��v0 ��(=
	���W'f6XB��	T�*�S�`� ���h�F�i�K-�]:�;��X\dt��O�c�͡%�wP�&iP���A�h� �z�9��h��v�8��#��ޒ������b�dL����U���5:2b��0��XaTe�ټ�IP I���;��H�T���l^U~/�c����G�����{㶥m�z�-]cŧm�<1�(El�K���J\J�b dG�;kv吱ɛ��,�,f7�|��A�H�N�<�ͥ"�茐��:�[X?�ԍ���#�o�$�*.a8Զ<��@���<�\� p�D��v��d�r�E4�츜��U�c� ,w���΃5��+��5�D�Y�{�n�G�j֐H�gˠ��~r�۳�^����ފ�߉t��3֎݄���5f=k���.Sk'm^�DM^��7[|6�x܅�
SK\{.YŽ��Z�腮��A�O��*�+������i_=�Asb`������[����P]a%���k���L��g	i���A��w?ղ}��_�>��؝i�Q��_β`'�B �1�!a��[�x�t�+�����p)#
@$���=@ٛL���A���>
�1�L5$����eD9$>3�~Msr
i��Wl��ϋ�����=$�E�7q�����2Cn5�LPм4���o:��{|��)��&o!���r��=x�Ju��~��¢J8���b�_�����pW+����BL�l�h3���q�c��Q*�࿺��.���ڥ"����z��=r閱��>��>�o�4|�m�|��ycI�B��;+	�|���#��m���4D�q؀��TSh���\��=�|��Y���t�:�f�"���̚��΁=[���^/�MA������v�F�E�2�?�c%��K�R��Qu\F����a�&G|��p,��D�(ͫ���B��2iM���F~f�B�х Jf�jJ#����5��zzfcof���6���;^�#Z�7��4ɻx� ���z�MjB+�BxŴ���`1���b�ߒ��W�}���6�nVZ�G���x����z:���X�mY����(ܺc��h�z�Q��]W	јEC&)\�Q�(�Z����]�g���lO��X��)�@�����6j���=�'���SB�:��V���6�`Ծ��$��tem����a#r�ڟ�$a�]����%�>�@r�1]Z�?ǥ�!r�ckV�K�X����$]h���%�_Gk"a���$�_5~G�������Tl'�\ �b�~�B0�^*�*,�P%�����c�.}��=��H�ܙ����BG����7T�7�ݗ���,��V��[���׾G�&�Tu�KW��	�4�4��Y ��N��1a��N^��+ɣq��ܝ� S'o��C�w�n[��$F�����_f���)o��f$pC�V6��>7<� Vq����(4yc,RNv>�[�_����"��������[y,� �K�mFUm��}���X���zd��B��B垤�w!%������7��/W�P�9��@�N_>_���?�=�t-� � 0%��|�5'c`�ˡ�8:��^b.��j�mc�#Ed�OP�2��������"U�_��^�A
I7�*'g/��ڪg�Ń['&v��j�c���QYi��ߠ��f��I;��
.A�@���'hA�R��]�p�[K��@b�r�W,�ۿ��ʌ� �Y���ROv�D��D���@����+����u,L�{�;v���ֈ�*XnȄ�e`����Ϟt���a���� �:�ޫO��b�ޭ�k�5�=�~�#ŖT�I/��]���/�?� m?�"�< �JDV���l�iJ��W������<�Qn�t�$�o���	��_��A!��>�V�`��J� ��Z&:���k�-,~شt���4����y�ҕ�=�wE���%$9GY⎜U�:?x}��/�p�8��	_��s��k����[��e�;F  ��S�J	
�^��������4�-f}�\~��-�JK���$��5�� �@����,W�`e�C�+�m%}�1hD�9��MXChj����C�O��t��&�y���l�G`���tP�F�to��,!IG�V�<ʆR�T?�^=}Y�=��OX�r�e��f�c����}^²p����˲L��v�4v�_ 8��X������~��7;�D$� S�������0 (ۍB��]s1bΔ�����?*qD
���K���7'�G�{6P�օ=��D��DC4B��dBwxǽbgw����s1#{c�}~/y9D ����*(�'�t�ȭ��|W"	X� �_�ڗ��N��e����R���F}�����ʦ��HeEL��������y)k~���X�����%Hn_W����Fc)����¾鯵M����A��W4�Z�Z� �kH.�֭Z(��o�9Hr���Oc"F<ǝ&��F�tn2�n�%�ָ.Vi�%1A��I.�3���a�`ȳ�g:���
o�D=͝DYQ����N
��9 y{�+3��%"{9�����f�1�g��tL��ꕼ����"�0�n��V��������3q�!	r����!�%ah��"S�\����O��ڷ���fz���쭲��򌃜�R�Aᤨ�K;¿��կ1^M��R!|����L{0��=p;�AR��	���$�H�} � ���{ă��n$q��K*ǂX+���y�����i��z����l�Ҫ��$���sm�Ǜt��/�w�
�ֿ��@I�_�_4�dL/�U���̓m��oO�ڝ�[�ziz"<��]^�3f�ԬQ1��k��,�l�%���Nq���
㢽���:ꀈcˣ�i%T����z�֐����,�Q%�b4פ����C�I
#�h�G����3Mf��rO�"����NcΉ�zQr��qڀ�u�� ix/��s�
9��
�y���K ��=4�&�^T���3���1,��ű�|�5�~���iv���,�����w>��F�χ�^��/�Q!L���ѐb�ez�Q�"�BtQ�ʲ�j�\��q���g�ڟ$R�
6FKbj7��a;���>^mыPE~�v���ĥ#�T����>ܛ�0NK �	�Ko�܉�k�"j3J��$k�0�4>��A%���8}�G��:���5~m�S��y�a}���ϫ⺁����r P�����Ę0�M%��ا�G��2�b3r
�!��7�b��A*1Jg]
����GՔ�t
��1�Fa^�,}C\j�(#
�~�3.waIM˹�f���!N���k#V*�#{K��)���hr�r�>z�ɉdU�<�>ih�q���i�,���n8�&'Hw=TA�Q��jm5���$�r��S�u,�

'��H��E���iNc�O<--�����0M����*���ʃ���<���p�;��h]�d��ke3P�ocW�g�����_�Y��"�Y�J";��An,'�96� �)���I�[HdF?7:�࢙�#@�l��-�~��5���c��C'�KXPE%�833B���G��4� H��h����&�4{h���F�p����d���V���Ji�Q �_��9�-�d%DyD�o8⭣�K+M���8��U̐}�0��QL�݂.]dRM� & u�{B���?�Vp�cJ�E�~Um�8�.����Ǉ����Ĳ���Xz>v���k�k�@�[@����;x]���$�ZS\�X&t�j&^X׎�=�%�[���x��1�	�F8ށ9۫ ���Pk��^������t�"N�W���ٟruxm�7��J�,Z$UGA�\MHB$�Y)o��#�S��'َq�}��+�S���7�CٻV>�7"�>�/�u'�k1D�q�/N@�Οk�|�	��yT((�j'�������.?�#l�����KVۧ��]��4�a����'X^��R�������{�{./H��:htJI>
���m	���|8�^���l�d�ԏ�$���G���HKQ[��ur�.�����A=�X���J�8�y+��sv(�&%�؇z�"�=3�o��:��Y��~�Y�S^��f'��4�!mĊAFO��Ɋ����a���{��NhH�VR��6;d*�����0���1�kCٽ2���p�#���ю��w����2�vvZj�"�:���]k)�̇1����Ji< v»Wor������ϐ��<�̇�x� ���} MY7`��4b�ZC#<!�	
�}�����hY�7�����kک-���u0�_O8�eX�&))OG��O����l��ޑY�>��
����Q���e�\�p�E8s�e\��#�(a�&ou�T�i��e�U,D���u�Oa�<�h~�692#M�J�E��5)�G�M>��V�6��E�=4�=�nc���S�2�*�yu����	�l��fα��J�U>l��׈c�+�]�{�s�yg��q�(�_�6�%�K��$�ޗ�����K��?�S�/����y��<.3���*\�j3:<������ayV�:���f�?���V[Ҥ4��¾HtÑ���q��p<�2 3��Da�e4�S��X��mW���)�����-�ʑ�Q��;K#v3�y"�/G,^֬�$ng��v����#6z�6+�ma�;��G!��D�lU��k�)��mZ���hbEe0�G�}����K������}���2r���v�[=�6~���Pb���{�B�plCw&�<'�����L�.���ߺ���5�Z[�jJ�KO��@��A9	73��kt�2o6�+Ǌf�rVcs���_yꋭ�z�Մ��G-RQ������,Qzި����vC���b2hg��g�U�F�׼J1X�h=u�,cJ�4���0��a�0[8a��G�[1�?	$��PL2�����7�8���n׽@M���^���ޜ��zx:��H�"I��$?>M�>Y�|S����2�*����!)]�
M�o�^lF�.�,�_Q�0g3j������N���S�h�����Q�P�� D��;��#e��)�AyU}��:R?y�T���I%�h���F��E��:ߗ�I.���k�w)�F[aj��$�R�L+��)��/2l�Ԥ�o̼M�#:��͂��qF�?v���6�mJ�N�=��v�`0�����;�"S��#�t�8x2 ��ɘ?�F)�Z�B���������4@�HtG���Pr�C�RX��k?t��v��#Q�}�d���
	x[@#�f�/��&�D��u��z�U��f�h��#HZi��=S_LY%�X���$,���p�}=�̬�@.R5,��Q�s��q*\Z%��f������{��4����ʸ���:02�??P��%�˞���/'�D_H������5M��;���?uѩ�<����B��;PT�z�ϨbpFp$	���P�"L	��b��5@!_�5�k�Ӫ�h�k�Tt��¹���yG�4��
:5Ԧ�U�nw=7m�u/M~�R��$M�>��[t�v�΅�w�-�f=S��������,±NY1��z���+����$	0�_le�����=����qX�*�b����L#�u�I� T@
kQ�n��I��?��.mٖ����Ccd���J����E��W��/�"w�a[�0�o����rj:�T`X���G��*a�%Y��
�mdB�X"So<\�=q3��eȯ`H����^�g�	1����r�j���O\��'e��P�F������[/���칓I�|�O�e��ʀL��:�������V�?Fm��'�l�bt��Ж�C��zA�)����R�5q���	x?�f��5�'�}�K������E0(�A���7��=��I��<�%�U���L�+���r�nr�m�!-s� k��!��x��������n�FF��^���T��� y��^�?�~fUό2	�P��B?B��e��*0��
��cI������K9�r�\�{<ݱ����ü���<�WYn$��nJ�AI�;D�l^Sk+����Z_>�LKt�α7�!ݵ0!����a���d�F��X�d��nnF�����y�q��i���5ǥ�ڽ}lS����]���0�D�t� ����KgQ�	�H^j�ߗ��=w��p��Й!i����	<��'���?����T�s�QY��+�v�Z�e�:(N���L4��D��������{7ŁvEo��qo3�=�IZ&'��0����ś7�����
v���%$��{��ӂ�y�!ȃ��xp��y�A�,�u�����d'�r��SD:`��2S����/� �ܨ��`m)�z_�ӻd��A»e0���P��9���C�Y�I�4�P���{2M�?%q<`����wkKsPX�� ��`f��H�冑7(�aG@�Fp�bB{(���*�c�]���$��Y��vg�׷b��b�Z����K�uOB��eD�. ������ޠ2|������)�m��gC��O�z�[l���6s��nR�<�b�����Q�`�@�"�,������ȅ^�)H��\��<}���/��(����]�җV}�ӰE:Ya*�;s��a��Q���X�
π��eu7]f�[�>�s_��~1�N�i7t�O_��o�1gܢ ����U�R_g�:=$o�_�y�[\vvT#=Gi���+K�����mU��^'���
��?��~P!-��h�&�b��7(ߌU�'��w˥�� �o!j.b�})�c�j�!v�=�s��o�� ����NkaK��Aó|ݡ��bI6��%A�[q!�#Q�9�(3�n�`�Tߞ�d��3A�u��=}�a�K����+���mXpk�0kо�^��R�I�5��W<��; S[.�Q�z� ,����{�-ڽko��%\,�h_w�S��&lz��Q���?��Z�����6��ٰc����0^k��������ծ���t@MK���~j,�vq�b��������/\���Za%���3U��L����V����~{G���ZI\ n}
(��A�{�Fd�F�x!P��*�J��\9W�=/w��Q��4��yT�쫰N��A:|��
w�Z�V��:�kuNO���{q��r���pT8p)E�� �߃����İK�S5"��̻��؛���<9��L�B»����nWJ�c]�Cwdc�g��}Q�iA����k3Pqg7e6��>+N���gf�8E)C?h���DGV/���[c�ƿO�\R��(L�}ҁ����	�F�$-�M!�����<�"��#��LP0��g+�&[`J����&��:,T�q>��\ۅkmY] x��,��	 ���l�O�bL�꡶|�G�/�)@��=E���gmڟ�@BG�$�^���C�#�mz)�=W/�P:ݮs�K���Nϗ7�k`ͱ�9
��$����UHRh���x|�})U�-�q!�L��U���A��������8�1=��L�7���X��7w�>߁��=�j
Q��4����c���>�6�ۼU>���D�|�[�8�p9͒�J�Ra�� X' ���t�_mV9����HX0��fW7�@�v2xM��C�	pǇ
H`>��4r�K"c�B-ȶ����S��)�"�O԰��d�5�AKMի����ߌp'	쐒G���C~��u甪Ȭ��V! �I���=g�+��.�q�M�i��������(!�$�XlxVHYEB    4f62     b50C�"��yڛ� ����u���-�s=����l��V�ULP��
d܆��,�--�,����qoZ��2R�j#0��Ҁ�$:I3�\�^'"�$�hw$�mlЃL���b�](�-���#i{�0o�I������������ԭO&@t�x5ġW��B�줜(ݕ1�G��l@Mӏ鑍b��9�7/��Yb�w��+<):lۢ���т���%��2��Z��ů�B�Ϛ�,+=)g���w~1�0�l�&���훥�<d.9n�n����m<`ԓޢΕ
�M���la��+R���{X�Hf��CS�c���\��DÊ޺�v`�,��ܽ�#P�m���/eZ�M�������	#���� ��\���O��;G(Z�qH��!�ǈ*iz.4�G��/@R�v�E��Y1�S���~	�Mu�QխR��8��v�cZ�B|� �Ė�=��J�j��.�7�Ǭ$�4� o(D\�<�R>C�Pd����*�vE�i����U�DRPb\�.G���%�qs�}^%���s�aZ=i��D�d���?�!�r�I��I��Lb0�c:ϭ ���iR�W	oO����{���ۤ���?%�*��Ґ1';��uO/�U_�:3���#]7�d��Fn��+��E�"��W�����F�F籕�u-�yJ�MM��*+|@�F��D��@��p7|m�[w��c�W��8��}���X������5/��g����N+
��Q߶�����C[N�q���f߅�����x �l�V���+��*�|'@ᔏ�|�w'nd��`w�����M��p����`�!�������n)�$�5z6otk��5X}A:�>����7�Ml(�x����!B�e�b�����!�VǕ��bH3�X�_�H���_z�g��ѷ��ϟ����OR�q�𶛶�ڷ����ez1p����Z
˕_�=2i�s�~�DH�X =���~��q �/Il�<�Q2d�h��X����A5<@�:>.�+*�r�E��r�ō��&[�L`�G�'�0\�G�Z�cb�ifĈ$a��^HT�+Ph�����=f��ɻ��|Ք$�Mx	8�ag}|���Jp�d��1"��s]�S9���HB�bA@{][�wbpa��K�����>G<v��4���d�>�P߻$&2K�Y��T7Z��_�[R�h�Ί-0z��* CrN}[�pi�Q�^�H���6�r��z7����8.=n�w�;��ξ㒈��H-'�:���~��d��,Y�ʃl���
�7Eyo2�)!�4M����/b3�ei˶���ÛuH������Ӈ�7������$�8�0�����01ܞ����i�l�v� j6y\'�������`����D[������(yK����	�c&pm�!�w�buւ�V ۑe<6��P֓�����Tƅ����R|�@��@4�1�-�Z`�4�ެ�y�j�lX��<�0I�U���w��C������ώ2l�v2�މ��صT��`��C׵z�Eԕ�'%F�^��v�F���յ�T'�DK�eXL�{Α�W�9��.��zF,~�`fH��{����T��ի����w�u،�hiQ/�seX�Ow����PgAм!D��/d&������Ք$ �Q���������$7�'(u��X���zTk#g�ڥ}��G���fj�0ǈ�s\��|8���hxG�����N UIʚO�GK\���
̭�썛��";��A��2���뙹9���n��򩋊���Z�&���Jj�*8s�u���S�k!���8=b�L&6~�,�%X��5��,�t��}>�:�{4��c�"�7�oc�htU$֡U�]�+Y�H̪4��g<���ߧ�Ql�����+#���ʢ�W0���tl��+���ӫ�L\욢�-w�_`�B�����?�Y|���bT�� (Èݨ�R����Ù<-�y=�B��GĄ��������%���B6V�kE%�mZ��#i1�no�&����p���jߏ�z%��@����?�2T���b2�H>V��0��x�-��d_��vc�6�
1�����[��+�9�2j%#P�L���p�L�b�e7d9	�Lw:7�)������)��gѹtz���'R��LXrZtQ����p���rw��T���|a�����4�!}�y�\ʳ�j��p�Wǟ��-�����LdH�\��5!�l&43W�H|_ZoH�i�>J�J'��Q�-�C��� e�L#X����ϥ�|¡R�h|�=�{��e|�M!67�j�1u����D��NI���x������/]�>@�#��Z��.H/�PƼ/l�Ugy�1�f�o��3R?�h�Jz�qv}���C�����nD������j�#)%��:4�f�K�Z'�:;B/��%�W2<(�s;!� ���*���ᒑf �3�1�%��a��آ�v��i
]%�D�XD\��Y��Py�L=Os�X뇉r+��\����H)= ����<MS��5�9�dU'W�*�\����&f~������P�QɰW�y���6Z�k}�':��P]�{#~ʢ-�]?���=�����DUd��*�#�WU��:��J4C��:���GęWx(��`0�����0w��HX�߈W���+u�q��x# ��d�f9.�>��1[�d͖�_��T󢲰;���x��c�σ����6�ll��k7���b%_�mjx�4cX�Wp�෸(�hҿc'�n6��W�Vt�����+�b�!vS*7L��Ӗ@>�ɾ[��X���ki��^'U�b�S_V$�6�̚w0~0T�\�T�J�0��oIӘ"	�Lw��O%�0�͇����}�X�.?˳��=��`��Iҧ