XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����&����^��(L'��c��S��)o�7d����G�u,Gʊ�O��Ð��NTC&�/���>��Gb�-u����m�k��ȣ[����0�x|��2C`˾#fOo�ޠ�X:���3Q:��a�"�
w�mC#�w �-�>����SL'�gw͜f���C�?2����%�P��M��=��B��^�{d-��ܛ������\=J��eڼ�U�@��@I@0�n$�=X�]�kr���9� _��-|�0�(q��� ��\g�cY�(~ʵ�a���"B���<{�~�i���R��Q��ˬi:*��qv���IGo䜭t����,Gr�Ե�%�'��sXi/�f�|����dݤ���o�)�Л� �aU5�!� %�[�;?#�83)��#�px @�`�q#�%UiYBg�w+�8>�:#m|m�{~g6Y�tF��N�	��3H�Ępl�J��-Gt��f[�#�|x�K��^�#��fg,qQZ;���`'�օ�~������%[�b�6�N~i�t��lDQCN�FpAA���%�`wE�#�q��*`{;��X�|1�F�?!���Z�NX_�%{
��vo�F5vem�b���<[�56`=B#�*v�\����΀m<��-SHI<hlɼ�T@���'�p�R*�>j�����m��jJ��s��{�{o�a��N?�vӻ��S���(�!A�>�O���<<��4�����=<ɤj�]�e�*
�ϝT��n&�_�*�4C��=���Ja�h<�(CHs�b�L�	��M��>�XlxVHYEB    3fdc    1160��
aǝ����J�
�Ǡ~3�p�j�����Z�o�}},��r�59�)gc2����0HG�XM:�6��XV�o�N((� ��}3ڄ��{��.CQ�(� "Ȱ�&�%A��0�F� �|�Jk�f4��"pwĺ�g������0��"��tu����2�����2�g���z�?9|p��K���;��u�rg]�G
��Y���c�Dp�ǒX^L3s�Ę�!�Z���<Gg�+�q�]t�B�45"o��ˤ���l���z�§/G�#fz���.�:(��5�dȹ�w⛎�G���+"�5,T�C�V7��Z����4��j��94	6��E����˙�)��]`O�~�$�.fw���^?*{�Wd�2L���؋Y+<}/sOH���_JA Z#8�Y� g��>E<�o`�:T��7�5Ƴu-0��`�_��0uS��.�����B�ʱ|�@/�y��ƞ[��wY�D�ak_�в����YrHo�F� ���h�m*��}-��.Jc��o��&h�e����$ ��腌&nq�p�	��Kl�	r�?��4��xS�w�,����;����?�dp��@_��9B�]�ƒ�k�ृ��r��o����S�9��4`��j�8Fֺ?��Y�!��ѥ-Q�3��P9�!�D:|B�i�mJ�)��9p���=����i��E���*�Q�����l�K�(������*�F����@���9?��
��y���" ��Kf'��67@X >�f&�*L2M��
pH�	��B����:/��fa���#n�
�鮫5���\L�.�����x��׵\���]bϊM��Q4�/v�&�����w�0230ϼ�\fL7�j��
�ǎ��7d�|�q�g��O���H�բ��
Q�D��1�K�U��Zsvw��i���kQ%������[��SU�q@q�u��O�%+a��ᵫ,���U�wh��q�iZ(ɏ��݉q�ks��w��O6��\�Q���f�_��͢�6�}E����� i0~��������w�s>����ˈA/��B���LZ�,�n��3�m�%m��6�y���-�^�~T��7���Mh��	b1[ͼQ�N�1t
���8<��b��	�{��DK�J��ښҤ��EB�~����s&�3ɱ��X���z�E��a�C�t�_;�떕��������]Q
}��ɳ����� ��<&����8P;d!(�ׇpg��k�ow�ۛ��um��ZU�+�Ҡ���4䴯dۀ�A� ʤ@s�����n$o������C���?w��~���s���F�c��O�|�_b�3����d44#�k�4�mU�hy$E$;oT��L����x�X���
˱P�������p	N�>�o�DD[��PasMZ�-���5Rк|Ԉl��\��W:ӷ}��lH_��5�K"9���5)���1݀�]%��ؑ����EտV��~�!с�L`�Ow�H:�׻�tϱ{���2�d]���!��u͠
	���oб�D%V�A�0�Va�LK(��D��.|i��c΄��N%}�|�q[�=��YK6�vD��Q|�q9�@��2�D �c���V1�+�gav��Y����=���MD��_����Hv\
�i�{tפ��	SI"p����E�Z;`��O��<x7ԥ�����������Su�I(�Y��0d�'���[6���TW�*�U��Y��C:�GP�+�;�d���A3�k�)�7c"�ӻ�p&,�i�%�uu��G���CDJF��z64!\�%�r4�]���ܠOI�iQEc�/߄���^��zw��/Ox�����=����Ȅ��=Y����������_�AD�����S��/kQ]�ܳ�2����F�$�.<�K8RAYg];��|�!$����gES�EMi�nJ���v��+��"8h�Ӊ:�o�w���J�82�W�C>�,w\3�[� �s�z7�1����S���#@Q�o��In��%��}�s�����s�h��D 5R�{�ק�8-���y��?~���i��1�����)���)Q�C����G~Kq��(6	�5�GXtÆf�Ԯa%�X��/���㺳i�;��\��'���н#5�&w��`(��!K���fץ�j��0�T��y��R&]N�����b�0�q
Eg�����(p�EM���l��u{Ge��ҌҐ���Y��;'ݿz"�Ģw-�Y7�����%t��b'��fw;�x]�ʳB��BWr��y�- P^B�h��o�5����6`v�f4�A�_	N��p'L6#8�۹S��@���O^�F�uեx���.�W�<�?�ө*���q\ۻ����V&:݆�}M�LX��Nz�>4�G�m�a�+����H�n��e��m;�,:�����(�"�+�������ۘ{�%&=^<�(>��?��)�#:� P\����)�����/<KL��l`"�Ǟ@�![1�Q�!d�:�ywk�:N��I��߰�b���aK�I�7B�D}a��b'�P��[��]R~���ꅿ|��91�w����	_��o&��`��I+�Ȱ`B�絝c�v��I��ƍ^�|J��t����p:�]?���M��-�\�`����o�*'�=�֑�~=C��f���oˬ./�!�����%�pI@M��t�����y}5�p%}�߁�B���d�,��!�yJ6v�%7?���C�z�I��1���>�d)�����5���Ua��d��4��0ރ�|z^��C~�a��Ovym�M��.Vx��&V��=��8E��%� ]iMa���%Y���}��5n�z�^Q_�ݭ�8�����2wʕ�4Y�I��q��A���N~�>j|h|�A�@��'M�X/N���Xǐ�"������F��Swf�Z�Vӷ�̏�:\�c��:Ӳ�Z��쏫b��X�`�5�F�/
L���ͻf\��څ(�s��]�{���p��L̦xC����)J��}������&q�<C|C0���Ғnͬ{��)����*�`�������
���\)Dc�����*�˲ʱ����'8���o�w�t�=��yM�~�Y����*��_������l�|x���<�`��� ��P})��?��ݷ�L�~0dD��ы X,5s���f5�`��~	�&o�\1�}?��QN0!��i��C��]���v����G	Zp��L�dU�
3�c�X��r�*X�އ��C[��iE���D��HN�"��B`��1���lB9�$��G��8�TB~ C&��Z��f�'fd��PK����հ���Ŕ�c��w�o�ُiwkW�,�t��}֫~C�kTj�͜�޻�?��D�5�6����j#L��%S�C���kyBL�S,F�-3i�%�_�〚G?0� <��!nT�MU}��L��HTbK/��v	exewJ8�+7��/7��K�xoou87{e��ܻ�W�hy�Ȱ��������s�Ɖ��=|����{m叁`�/�(~��0�֑h�!��,��s���S]������N˟`�����t��J�nv��B{��x��cj���zL�rWٚ=�Q!C� ���zT8��p�{1W�)=��������p �%�}K4l�.�XL�h����)c����我)h�nus-�?,Q&���u+W��(k�d�X����5c���	-�*�(3bO0R�[�Q���c0�	��x��^ �ăIyz7:dTݦ����ؤ�^�ԙ���]3�f�݆�bՠiq!=+����!	2-�~�@#�/�ׄ��k����ߙ�ִ���W`��k�M��=1�|�	"`��ʃ�=���;g99x��8Rr��{'�\P��pYT,�|�s�gO���M�Ɩ���N�c�kX�)�����޴�0�iŢ��Ǹ��h�Я�|���LI�wt3�>w�4�\Qq/n� �,�}�i�s�D��ˇJ�#�A�-�T4���_�0u�7o_�/c������-V߰����	��F���,���ܞ�NvQ���n�5l(?�^��B�G!� &8�Jk2FJ��kJ�aL�j%W}/��QT�T$#_[��Z�v�hz�S�=a���o�:n��Ӹq@o`s�L�D����$9\������,k3q�Z���~�e)HZ@�4l�@87�?V��+h$M� �􎳚�YI3��
���Q~�-�*�mѡt���A��\D_�i��(��]�aK��8c{�2�|��?P/�	L �s����{��XN���r���"�3��#eI�g��9��3 čN�!�̕� 1�l�h���AǛ�F�JX"��E�MDd�A�N��̊\gė�?M���e��{�0Qn	M4