XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��FG�ʙFZ\Ѳ�ѿxտrc�����G�O��dn܁��Pl���]%Kv|�����«M���V�r՚ �*�bl�+a��X��M�F���rC0j� <Q)��	�g�.s?�s��l���,3O��w*�5	5�˃kCk�
�F)�y��	0�2�ϣo\V�7��3F��M�w���=Pّ$D�������Y��<���NS���%;�h#�+\4d�@���3�?,mNe��^��Z:<�n�%ɬa�$��	`��t���BV�??���q�i^\1mŪ0f9vܫa��13� |�%v��@�Dy.�r�b&j��<�=����;�r
m�C q0�9'6ߒ��s#�r)�|�k������V�Э�3�u}K���� �&�1�FG���b3Gs�:s����w<�pSjb�S?U-i_������e��~)��ⱔXu�%mshD�J��te�w�tA����9	���$ݐ+��/JTY���_4����o����55*Q�D ���'�O�N�(����{_h�¿��,�PSl��X��I�S�0	�9F�� 0�{���ϑT�a�ʷ�q1ȶ~�*���?� ��b��Qf� �؛������@�j%|�ђ��f6������bC��_q��X�ƭer�@��<h'���*ɒ'�Gq���j�c�+����`^�zI�$l�7�%[���LPK�(���F�*����A�4�BmTBt3h�<G9�N3�䡻�EI�6U��=,�261�XlxVHYEB    1a2e     8b07������;�I`N,��BAz":���7�E�1���Rh��.�-����ؾ=��I>�w�K��m\+��.�]�����ߨ�X���1(@�Oe�/�(α&<�A&kzh���/��o/��;l{�x�� ��m���h������f��$��:5k�.̵�����*2,s��e6�^a�����~k8�I����0ՋhyC4�����G嗺����8-��y��L`\wq+���ɛ���W�!��hu��W��$+ A�OLg����m(�ޭ�U��	'�/�����åO�#6-pt��<:ؙX�����D�
�7�b
&`���,c��`�KP��L;f6��0�H겒�\F2�`������I�S2��dD�(�h! s�v�t'�H���t����ſ
x��c}��d�^K~p"m+��_F�q)�hj�q��C�.�I�:"u��)ءߤ�9�܋Թ�*���߲�1`�Yը�K}4t:c���3��*�+hD���(�lf72 � ����_KA����!�,������ 
�����Ⱥ�@��&�����KSips͎�f�_X�s8��`@J�]_luK.��٪'�}:��b�Y�ӰM�d��F���^����tvݛP�I*-([x�1�������}H���y�1�ժE��fS`�2إ_l��`���S�A�K\�/�@Q� j4q����y���AA#>��jx�����P�f�՝�E�M��}��ƙ:��c:�A{m�u���;�&��������B��Rh�Y��È{��!�HxM :hg�&�-ׁ`�U�\c����`�G9@G@�\�GnT���WW�ҳO��<CK ���g��0���L���Y����m��Wuзg�#��˗�5�eE~N�l5K������,���ǹ�<�G��d]�0�0(T����t0�m W�p�28C���4K�!����}�Sn�������f W-��<b~�s�qO���p���~�0c���� �y?:$z��/c��u;0pe~-�򡓄�E�OiЋ8���k����b»��<1��I}�dG�3 �URY:�]
�%�?!������+C���fUI2+m���q��7ǔrb�>��:J)@+Ўg�:�����Ȁ�WE6iG�h�2�t:�*�5� ��6[��$	�(~�"8��Ā`!�Ug!&�B*h6tH����`�p�%�g�� �0��t�Q��O�:�b��Sұ剱��B��b]�w�Ũ)l���'�5������'KL�2�Up6DJ�yWeus4��p%�����:���ONg�P�w+���>�35X���s��xf!P��Y7nrq}ձ���b.��N�{c��U��b;�9���KƑ��	�i%K92W�T��L�?��:c�I�����R��LL#L��, "����Em�
yz�Ӗz11��(�3��6����K�Us��g����'�g���vOmJ��Ccm��K��-;�� ��JrSX���U��6�莶��"g��z�%�Qq&�b��n������P�!+�䗨F{]2rL���fq�U2��+��x�-,7�j�xJ҈	�'��D�G�ɺp�_�$^$�}�N�߰�Jp����H7�A*��&�~�`؜�[B�k�:�ak���E�
Ii�
4����e1Q��^@��4_:�2~Xx�P{�bt��bሤ�h�|-��0��Z۱nֹ1�#*"��l``�$��g�ϩ)���L��]�đy�;hg�L�z8`���@Ӈi+q���~+�Xާ�˶�����(���b�G?�����Jxee�Bk�#�PV�nS-m,OHw�'�����i�ou�*����+�T��cO;���GB����v�M�[�1�񈉥j���=��c-?fn�A��T�o�3�*-����1�ǨN7Sb֣$�߯E����|�V�������N	����So�As��̂I%��p�RW�ε��������;��O�E���Bz�\6��g�f|��Q�&�П��0o��}�kK���X���Gn$c���/V)��ɑ���Sl��D$ư\gm:�d�����Mn��&s�XS��ig=�ñd�.�L�{��]�#μձ�c��/��*e߈���o���}�����5[к����ђU
��Q-6�C!����f���qA���kԎ.X:x;