XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P�<C\Ţ/,jn�q�n32:����k�����HѾ�Ъ	,�w8~S,���iK��O=���C@<�*x����`O ��l�|��7��8,��s�K��#IY{��Mp���K�=�]�z�<�.�UH�M��q�ߦZ�'�崴+LqLmF!"v�6�X�ޑf���c�{�3�E�;�e�.�(��j�V/�+��E�K�1� ���<����
�3����Y�l����h(�m�L���7�~��)_\͉7���3<��X�jv���1��Z\���F��k����3S�D��Z ����GC�?��]�����S�#\q�L�jz8��m&�p���ۺ�O�t�f��u	o��*Wj�T�=��ث�8�a�I;�K�4~��'?_1�S�Ѹ��m>����7k2�tG�tP0�~B��\�^��ؕ!�C��oG�X��-h��2�F��$Vz�JM^lܬ(]�o�l���[1ûY��@<���QP|��`�=S+y�Cl����e9�����{���ha�?,�U�8v�4g�L�Y�[X��i���~˲�����yk����\=�})I���>�������,<z�=���Pᒇ$��RvdB+Ĵ	�?D��2+�hP�C��Y�<\�'xZ��_�<�]����x�L�և�k�||4ڊ��UP��$�:�|�Nj���t�lwQ��0�ᓜꬤ�SY�a�����^d��:kI�:=A�+D}�{����^�⩠��Wd��a��z���j�R��XlxVHYEB    5cad     f00��(��4VC��p����"и$�������m7�8�+Z�x�����XV�n�6f@ox�Y
�m�?c�DlCS�����7[H!̥椾���S�����N������d��Cσxռ�ݩ�����^V;��6�ц���=����
#��+���O�r�S�k90�,�p&�yw̯��4��h��<��8�}g	�i���/�Bu#b$��e �-�-���K¯]�8mЁg��QX�%�=��J�Y���{�Y�	{����|Ƒ'Uz/�ǯo@}�Hcg7�pW@�
L��3VH��f���i�=M����n��4����z���}F'�=��佫���v+l�G��Jc|��[������b;����n}��e����&
��6�n��I�:g������Q�]��7���;F�+��L�������*h�7�M`����U!��뿠8 jp��9K� 3��(~�J���i�����o�5��"��e�8pA�^?��n=�ȑR31������0��`"A)q�Ԛ��F���
�8�x;8���kL7���UU����])�@� 3�zE��p��2��$>�C�a<(o�&DG6�rO��{4 �`�$�u!��6B/ʁ���U�%�.�c8jD_�#h-���Fh�\n�����C8�U�I9�M���M0�tD~Cy���͘q��`|,(��A8��tY�9�y�B�,3�zva�*1V��!��v�tѯ[t)��G����L^}��	z�3�����-E=�
����N8,\G�K����խ-C��,� RJl�6��<���>������D��X���*uj�� )IW��"i'�>O�D��-�a `~N�"NcFi���Д�h���)��Nt<lI4q����f ��e��\2��[�uǃ����?*�XL�5M�=\���	����|k#=�N��tW�L ��D�k��4�xPU�"lM, a�=��AO��v�\�J}A�=B�}�-������R(�P�>u�\e�ꗚ�m����{���hů�~uъG���@��k��C�&��k�X� �� ��Î�~��÷���}ل�g�baw��L7ߚ����a���+j��Q�3�{��e�{�|)��cӷ�䈑�!�M�x�)x4YH{D�&�+�@l��S<�~�X���s���bf[���� _*Kcv���|S�' P��A�"�㯹����ݠoF��b�]�l�M�!*5-�a� ��
�[�� \�/h	��=]����a�q�BSd�	�C����/�;�"�ŝk5�t+�����	"��:��̘��J%���[��z��+řa��N�[r�0���g>�a;��'˂�����q<P>T��K/@]oW�h"<2 o�FX֞t��=/�oi_݇�Z��Xur�/}D�zc��tY ���V��E��6�9���'���d�ڀv�l� ��hqX6���F������
ĥ�CJ��O�r��m�Y��o�"���EKjٞmev����7#|���ӈ]�G
I~/�ԮOQњ��ը�ia���ƵTk>2���%�x����la��cl+6^���G�gP&ؔ�5���j�������;��������`E12��%SN���Ђ����x���o '�8E��Y�wՓ�U��x�Eձg�����v�.��?~����j��%q�#�dTr�5n���q:m��2�*E W�?��Sa8����*2[��ui��X��A�ME6�h�3��
6f����nf�՘\mw�g��|��7�f�k���ùs�K�<���t���;��2k�E�֊	VX�x��>2:����ӻݙX�{��m	���!ͭ@��N'%_�;K���J�?w�s#V~�����������7�D�üoJ���Ō쾠5V�������	��#'�ʹ.�"׉�u���,�sb�B3[���|�I[�� �zX�K=B�P�7����<Z;*􁵪,5|���%�S��-nP��=�F�0�O;Nl�㹈�����bB�GM�䩟�[ԁg�n�s�Db�nGP*MP��=Z���bmvĺGg�~_��.��
�.�Ę-�r��y�uC����w�4)C��#T昧G�1mPɛ���0P9M��y�)��2o�i�K[��Ӭ}���6f���'�y�2P:,]�qah���~���&���>Ԏ�z��I<S�.Ud�P��(t�?tQ�_)%6���N�Pu������� g��5A�t0՗,E������*��������T�����Y��=<��<	���N]b��ڸ��(�7�q�H�T{���}��L�f/D	��ث���*���?!�m�*�3L%~1�s��4�9���k��@� s��0�����*���V��M�K�W�k%.v��|ڡ�Y�7x)OX#�7N��q�t�n]��8Ȼ���dJ�����1ֈ�3���'��'�_��˓��-�u@����&�$6�e���!������G�Еtw����{��Tk4��}b��R�g������=�:�v����Q���"���ƫ�mw��&�0�o@Η�T��p��a	�n�3�����W4�D�Uj3P�뾞/�����-(��"RIT����H-d�(ؕ����,�y���#'u��izc~d�[^����lXz꧛w<��!�P��\�� �W��-^r�����Ւw�um��bR�/�D��Ctw�o#n�0�.�_�l[��vƧF��@LU�5
���q����ȹ?i���U	~�kLv^�/TF����N�C�]:��S���f�4H_ß��2޲ҥC
Nܖ-���$'~rBAM(54�O�7��a[�>���%�1ӔF��u����n�Ԋ9�7����$+�|������jl�H�>wm!��5���Zj��H9;I��TеE��Prؘ�b��-:���$��Nȑ���[�@o�m���������9��5����Q��X�D��t�N�Vd��}�C
Y�>�z��k *E�m��сhpρ�-l���Kl�J8���/���dw[�j��N4AI�7J.H�d�#)��H��G�˱<8f�4,q�jZQ/��R��cL��ŋD\�������9��B*̖�Y̓�.�~��h�}t� ��c�ۛ7ٛB0�����F
k\��b�1���("¢�%���5�Bu&�,}=��!���H�_Э�r*�~�t��y�y5	�Z����X�uO���C8���.�x'�+{�"%�k�B��?��kn�6�ހ��]��$B
�oF����j@1��7)����~����/����;���|i7�UL8M=��'�0)Ÿ�'�"�D�����W��r���%s�}0��y�L��䐴�y�Q"�CJ�-�ǒk�,D_� �M�����E�^���W��W���c���8�~IQ�&�'ݥH�J�hk�I-�7�A�⊅�{<�{wX�CUM����p��7R�Z+������w�%]���� Yk��`����y&0��A���)�Pou��Bk����Ӹ�ʕР�w�����mH����D�_l3=/&}<�{u��P>���l\��lj�=�zo�
���s���Zu�cR�nk��T5W	ɋ�K�Y�>+��7S��/s�����uD�j�*�Ϟ��]^@���0���5�rڅ6��Zf�LP�.�Aܤ�����0"!�u��cl���wf�X�Z�h�:��M�3?��p�W��R�o�"�+���G�@�+ӾD��/7X����dr۩+MQ$Ou��kjx�`b�3