XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����;����!i��s�a!��q��q��Mq~�l��m�����O|I[�ߠh�B����A�Wgȁg@�����r6�ve����*����+�=������H���|riqwc��s6���ю��얨b��(�ۍ Hu�21\���|c�Y���a���� �:2V�|�Y�ki$�e8��J<�\�B�%�<=Z�To�q��������s2{fj�>����"�`�`��\�	vaV����
ӹd&4芜�04+,��$�����s��2t�Z�|nĢ��'$r�Qy�0�����7���x��L��Cݐ����2zX0i]9�Ӹw鼀����u?u�^����g��Gu���=UО>�Ҟ�ڛ#�S��D߭�,$�6���zM��
���;r^�ŀ���ml�Qs�$y�j@a�����1g�@44A/�[Bh�b�/f:Ԩf_u^O��O8�Q�AXH���Z
	=��5+�	�R���$m�����<�ך��\Q�l5�4�����#�4#�@�vg�X���N�@݇9Ȓ����åQ�����1Q}8�u�`_#��oxN�����f��8��p2�sr۰��+	�O3�K��3~�C�{]�-�qT��Ȯ1)��oAZ��c��ǩ'E�`_��w�B�7!N�zO��w[�h���m��q��.��e�r�'�nӗ3�)R�x8*�/�>�t��]��*��~����T�O��56<�͸j�eb:�e����QD��o��EY����w��	�_XlxVHYEB    241a     ad0Ra�$M�T����+i�ۯl�8b9�z���[߹�U��:���;n�ˢ@�b�?8���s����YoF���Vm��T�*̧�"i�!>��R��k3���}&��~О�q�"�mM�\�b�?���h��x2f��.���3��|Vڱf%�&*�+3�ۆ�}��� Xz��Aol���Kj�~J5�C���@���c���ÛY^��ݣ��Ք>S;���h��Xwd��"���,��zЪ{mh��C-�V����A	z��V �\��<5���P�`�V�VǨܘ���l�k�۳��z|�V?'��������:x��˅1jv�p���J������B�[��a��N�8�l��&nC{,9~�����zB#��	
��WteE��e��L"aY�0��M���|d��-�����M����d�l�bnP�Ĝ��3>�0�z��f�2�6=��jP�|�����~��'�[=�7��[5���#�u�C%��E��3@����I�r"�o,�:�	� �oU3̹����jh.��>�q�}n�Ӧ�#}Xrq!�3K+�� ��.�])�(���hӻ�$�ae�Q�'IY���nf�iH��E���M�)��������RL�W�v��[J�?3wo�"'��M\����	Z�����`7մ�kI��6���A�y��d���7%��� 	P�L��o^Q���6�YZ��pHN�STk�����b��S��@!�� O브l�];����Lg�����S�����Z���ڒ��,��ʿr�M;�SN�U�+������	�ĪS�D���(d2�J�.�L��}AgXe�6cX�2��)�)����g/�����7a�XG
���\-VQ�IՒJv}��L����k���b|Պ��(�2C/�
F70h�OFf��L]"1-�Y��KS������~�~��d���w��.�8_�6i��2	ݜ��K�u�5�Zcl	��S�� �_`UG��i�&��<cu���ύLɗ^�	�gv�R(���9@ְ4-d/���KS���9�����>ͽ� 3�+ �P�_L�M 5u]NXc�g|��1�R�lP6�X��C|a����.�3�x͗��cR���ᎍ���^<`��vz����p�;]���#�I-�7��R1lh�pz[��&���DF;ǐe�<�4���ڡ�� $,���Q7�dI����8� C̤�sC�H7A�'�V��'3v^�������X����7�h~	���|٩�钥�������a�b{ųgZ����ñ��,�f�;��+��Q���]k��7'��wJ���H����ЇlE�|��x��H�%P��?�h��p�G�������t41[�M"����(m�K���`��2�ғ�_�I��g���W�+��#�%�n�'*\(��\�P l�H�-:p_���.�R�B����+|;t���9d������O�,��T����Sa�y�;��j�O���U!Pɺ�A��M܋&�?D�/3	����I�Q�E@���ܝ�Bya��t�J�L���n�0׹�IS�T���:F=Z��x��l��zp���=4d���[b��O���l8����3�i��e��R�{zFb*y�!��~�]\�㾠��W��L��Ipp_�ZE'�4����]����{U�ڹ[�k�'�L>�͞�:'�Q�,XZ�vǿ �TP��3A��H�PK�_�>� b�ql��?����7fuY�KeN��BǴ��Ѥ߆�3�^�/��n�@�������j>dôF�ze�T���g�6��ț	{F����=Idݔ��� Pu��޳���k�(>����� D5�b�#��y{����ڽ��M9"=�E*��7��h�N5K(�}��W��ǆ**���k�F���TC��,�msN�J�X�ym�0����N�_��`���7k|��j���~0F��?f�/�c�:x�q�}9B|��c�=��������Z�de!LOYE�,���◺�A]b/]a�s��	'z(����I�7� �~���?�{ �I�̴�h����%�C��S�1�O��Z�P�g(�Q;3�8hi�2�*-��S�{�m����o����r��2�B�,�v6�8 \�G�mh%�6v� ��2�.b����Um/ࡣ�����GצL��!�g�X@乫@��cr�Ӿ����'$��@�SĮ������ҽOb�Ki�J�&��#���;��oξ*]ǂ\���lZ��k�x�M�1Nk�1-�>�n�6%���=9�|3uI���	D�V��=+��·�wZJ=3�&��.���v'�u��5�}�YZ8	s��Ќ�f2����D�:����$���ٔ˽��.��(�Z�`�*������p6s������������c��a.hz��Ď�Y.by��z!à]�<��d�B��}��j�<*h2m���l�ˍ�as���������WH-�:5m�@OVs�-3������� F�5�q�
��� %�Zyg�T�f����3b!o}/Z�@0O?�X�!g���I�w��،�C�6��-x�����������w���;N��*b�S�DAS��[6pN���C�eI�jΙ�.S�ۜW�Wt�?�8
��@h�|����j뗘	�9���Q<���ct���� n�'�z��� q
%�J1�VWa�Q�J*&�l��;��-��}���