XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������h4b$����jd����{(V����vV��fpw��aܞ�F�5���L^��ϱ��wx-{�Y y�>��Hf��R�����_��^�S8�	�+�X�*o [�6D�ˁ#�Ӆ���N>Ш'�c$�o](z���o�6�1:��9��<��Z�pMKR�7����il��7�%�̉mQ'T�t�ӏU�!6����6M8�qm�j�OCi��m/=}>�n�ASG 5�odyp.��tC�ڜ:����i��H�n�� �6�d�6_}�_vRk�*̘s�\>���[T6��Oa HH�F��_���%{��tѬ�;��LCX��a*��*����,_������ժ�$=|?.SjBl�Y-���H^��m���+T�ﲷj��ʛ��3�_')/S
��v�:Á/�ĉ��ABʕ6?S�S&�Z�}'Q�.�!���r����3 ^0�cFoE�
�&^#C�0�i���㻛M]$ߝB(�D!�&��,�bT���� "N^A�=X'��8�P��R�:��)�P�	[�נ�b0ݡ]�%��2�;�K R5�iQ.Ѻ��&ø4^�Z��D�͙���ߧ�a\�}˻�Į:m-��B3���+���W�|�<	�����4�
�����a�3�&x趴��]�h�	�'�a�R,��;���ַ�,,W^B3��'k}�ޛ
���ʚ��/�����SYB����ڏ�=Vob�x�e��p��5��C��b�q����7���>XlxVHYEB    925c    1a60�Y�!Q�[��$ry���l�}�q�(AN}� kx��/�Y�P���hń�p�z��FO��B�� 3v�)���l�O?;K���i�$\a�ۭ���p��Ua"ݏ�����N'aR���+qj!�9ވ�h �"z[������6{&dN_]C"��RB��,�[�QȽ������2u�(���pCP=����Ǜ�j�rX������/�#?*Ya�#wB�J�{EaY���o���FG�4�
6�d�i��r#[`ߎ1�-\>���>�t�Ì�+����L���4V�=B�B�%���AF�l�[!j��'ȲU��Ű��t��"r����^�������ݭR3�>YW<Y��|����c�n?���L�?�n��b�g�n	����ܹ�3'�\*(���֖�Z���zE�ְ��Q���'����+!��ҟ��5�;JD�2����hqQc
�u��+��gU��=F���F�a�U	��ϭ���8������7��׾�w�e�30<e�4s�ocg��<z���N�Ηq�s��wy�`�_��ڸw��/8���m�<X4\�G����>QP)��gB�D�r^{Rw݇��ܲ�'hIS&�	,� ��?��#x˭E\B�@� +�;�x9 ᇆ[�Q�;������ΰE��� ��70��	�O,6d�����%�g�1��J@l/��T0C����;��֑=�kA�ae�L��u���̑��X�����]ota�?�ٙ<�Ws�(d4Ӏ����O2�
�Ѐ.�uL�P$�)ncrቢ�gjwt���sf� s�]R�E1���D[.����w�����:�:���!��t8r�r�ե��wSU�,ͬ�NK��9qh�w��L���Į����k���b�y$��D#&�^���T�yH�T��S�g^��V2fm�1��敊<�ϥ���Kh������of5��(��Jb�2��!��ۜ�����e8�f�(�,���dF�j�6�y�U1%���KJ>������U�Z��Uj��z��y��ڀ��w��mue�%�z�H0$d�"#�po5Ip��dLr('�C�?w�
UR���<8nh�PP��������_��.�� vG���hL�lnD^Ny?ř^��w�d����K�%��a�#���-@Vzň�wX#=w��Eҷ`�r��ZeHϒ���
��cJqw��[�!����N		z`����~���d�4	�DV�EHo_Q��ש>`Q'��n_uR�����(Wڻ{M��Oܷ���|��4!Ex!��#�_Ś����8��ZGDG�r��w�p��l���d��E&d}Ȟ�c����l
�y�������Z�8QP�vِl�3����?SHɣ�B�P�U-���d�U(Jk�3�MgL�¤2�� �ad�Ga���3�s6���I��i�{fW���jĮBD�3G3�vq����C���_�������)#�%W��}eh��?�.�kbxDj�ݫ7`���/�$�%�H� 46`�b���9L	eZ�T�����̡���߸��Y�{������������n-���8��b-��~|
|�	���°5��'F�x��7D�C@Yz������'�	��m��C	����`�m�餰݇�s�л�N�n퇐Ք����g����?�h���ռ�80�f\~��ǧƜ2���cB��̩��Z#�u��ͭ�鰨���rCӄC�4�q�3�iJ�B)�K��B��`K6�H�=������"y�
����Q�y������͕+#��U `|$�<�5��Ț�;>������^�tcY�;(}��K�P�VD���PR�n�7A��Z>:�T|S��H ����E�چ�Cz:����2��L��K|<�Rt)��7b7QG�F*׋s�י�#�%�����]�0����?
�vla
�o=���E0d�@9%/��,���ֱNv��N�'e�.���������!׹$�z�N͵@�e�;xi2��ֵj��qE��.���d�u��)��{�e�<zҟ�� 5�G�^�Ԩ �4Ɔ�st�G�-���?��m �����,p5t�y��zo0�R[(rV�[,�:?E��=ͩ�/ؙ��Ջ� <J7���r�-B��Tc Zبv����?�ۙk�oM�f3Dĕ�K��%��N��_k��&߰��<Qǟwx�b#��(��\��b>��N`67&���q���L~����{���ğfg��i���R2��z�o�6gO�zL=<�.��Ti�`)m^�%w\Y7�;�g�-����R�#��7c2)��6od'z!�\(�O�P�y���N$zᥧ>�/}Е�tp�rC�&�Ԕ7�K��p�xE�v�,+���9���7���3�0�i��h|��ˎ�z������^D τ��&�ԏ�뤱�ʹ�(rj����u����v�ҍ���b�dql8���������,E�gs��@�n� =�� �xr�NaЏ�F�h�l+�8�s�a]����G300�L �H������������\�c-c��W��D��LP�j_���;�O�ы�����I���T^Ƞv���SҠF�>�����$�����G)�n/�奟б6̇��?�|D�ZJ���Ş�/2-b����(�H�dgB��	ja���+���s�j��'L�iN{��I,�B3���7P���|��aERKu���W�p*Z8v��V�����.l���`��P�R��O�<� �n�	N�o�(��Q��M\J��vp�?=k�|� ��{up��{���C�*I3�!4X�x�~��w$�9���k%2�OwJ����կ��gU��â�,����IL�7'lȠ���T@ 6ѣw/W���g�gf�eO���ߪ��8v�ZO�p��m��׹t!�Z�J�|���fE�^��;^g��t�����*�7�#�|'�yz��R@أ��M̬4:��$�x��1oK%K"��v���/���������]�fQ%�Jw$��K;Ī��k��U�vϰ3BL����[
ؓ9�Un�%�
�9_8Ө_�]�V����?+�Q�X�,�2�,��JZ6*�[V��s]{�����-a'V�h�H��}&#��p��EfFuT�[&ϖ|�����9U�����wEl~�~,wY[�q}v@����1�)u�W������\�`1T<�MF��@���b�.?��I/���v'�v�M��4�aG@���Nҡ��b�%r���ސ�F"�YX�u���wm�޾�]�M�!J���vj�.ᄇr"��X�`n�̠�G`��_h�'��� [��t��r����@4�'�����k��@s��x)�s��N�+����>�����S���i���f0�}��Sp֠#�m5�ۡ�;�Is�E�aP��5OQA�	i�e��]�:dtޫ	"#���Kz��;u��uO@&�M�8�
1�x���12HU��O�[�����y�����H.pѯ�۩_�?��U��{a]ބG�g��fC�=���za������B��
�q��J�L&#=�՞K���B�;����E�3��?h���
�c"����?�w�W�[u�B᱕<׽�7A:h5�� �~����S�W�L���ӝ�ۯ��(�	�l8V��b\�#�"�*����P�sL�7��\e�f�G�H"�z��x�w]jJ���탵�.l���
��h�;�So*�ژxÙ8'b�x�U9�l��4���,���<sejs��u�A��"5�g�+�]ZV@�`�#���}�1X���AZ��HH��A�"��!֦;ΐߤ�R�Y�he��'>�LK��-y��5Ϋ������d.�P��\u�=�mHz���
*��+z���tJ>��M�Gf9�v�n�I�g ��So�Y�nJD����_���t���?OP���@[���!�}�u�-���t��.�Y:VJ�v���������*��Y�(*i=�p�U�(2i8aP��DD����j�M%�<��j�I:���h��D����JB���VT[�D��X/n��9d�
�"`�+��Qn���Ǉ��ptw�e��v���s��i�ӗ�F�P侢��a�¡ZATq���@��y����=�[!�Mӟo���rH,+V4��#�� �YO^t�1�p*��cUt��"z�t�j��#c3�������
�G�s$0ԪӜR�oRe�CS��f�t��p'�ۖ��e9��
��s<��`�B�01:�*�vg%س���L- �ly�}p�����ǎE��%�fSJ�shP�HpU;���T���'+���Y���0�;s1̟���sJ�z��0����Y4�fy����]�Hq�7�)��A�Fu�s�/�8�6/Gŷ	ٍ���Dn����&כ�s�oi�vѭd��3��z:�&����Ҽ0Z���C�b�O�)�nT�����:�;љ�ڢ��ρ3f�����D>�`���-_�B��UH)�вF:�?�X����Z��B;�g�1���`O����{+���$u��L����� �MD������GɷT��)a/�W�G��7���<@��¼QR�j�e9��L�춱�;�t ���)�R�I����l�ҨsQb�B~;(8#Z����m"�i�Ys��kX�d#H�A	#�q�.C���GT��� ��Թ�������v��(2f�j���ּ�%`>&G����[Eɒ�����k8�����JA��_W�țq^\��G�G'�~w�r����d��|h4����.�[�|�w{��������j��� �-6 8S �<uf��Z�|Ig�V��q}���g��H]'�ݤ��@;+u{�N��v�0�GD�tc&�z���2���E�a8�ӭg <�� ��15 �V��1Anj��鴑��l&~�Q<���XQ��
�zAbEfyA8�/���� B�V�5��é�z�����΍�ha�g�D٦�.ȑ�ggT�^L^v	;�Q(&����ט^�y����3��D�Be���"�����P���AA�jX��x��9k ���vkߓ!4�sso�
:��i�(GEMǝ{��&��׾d��&��ww��b���(v�h�f��6�S�B�Ȝ�9o�Qݳ���Dt��6B�bkN�d�_o0a۳��� �q�#S�XMB;�[�n8H4��"J������}�8Ʊi,��Ϩc'��N�lFa��wԡ��fT�I���A�/0�ǰ�#;�������FȘ���������2�����~X�rs%63,���䓤��O��	�$[@
v(�d. ������M�>/,�B��CX./
]�
*q��wZ<��M��Kd��*���O�lPR\Fx�*3\l9	�X&C&�W8d����+��β S� �\Q�)��hĐ�Db�C����X�*�Q��^�r���P�p.�k�gZ��OO��8�e��CLŲ�<��=�;Q�ҷ����f����j��tY2>e+#�&���Y|(%]�h�(��G57��Yߚu���i�ta��m���8pku��è�u�JF�G XN6~95��!���/3��e��1���}�V���*��l�ԑ���aO�ei
ZL�0���\�H��ó��~����?��䨒�⒐��������.�6k�-%�2�b[�ZM Q�1 Ԉs�盟`C��}��)<䫱�O�}�d�y|l2/���l2&�[�q�N�+��[�of��u��\:���T�B���i�4
j��	.�c~���]�B�DdsT��2+�|���&dE��2��N=v�?ם���+8�\��q���\��p�0���������J�V�]�g��Er>�����H"�,@*l���T:!��6(B3����^��A�znػ�nJ>K��:��Z F>;�'��z�Ip�U���$e�?a[I�f���b� 0uV�1�*Rp��`��A�c����'�	����^ü=�F�%/rM��R�x�^�d�#�C�j�\�)��e�_�tJ��I?;��A �aa��hx��~�h�V/f���
��f�I�X����� }z.&��I���fF�
��t�+5����[� hx�zW�_�f�>�'�b�Y8���,�iy\��ƈ�z�
�0	���^��f,��h�ND}���H�a�&��Űs��̬h�c`Y��C�n��=�4�x�|Y#R�ˑ�-��1�<=��R���DwP#����U��Ė0.c�hxe^�+k���ES����}s��Q��]V�^��f]�?�9Z�G�4�I�Wy���|�~�	��lՏO�u��J`�){���B�xѰjo�deQ��-iq�c�\Q3��=�_+zh���NAd:�RU������:V�z�%P	⡝k{B4e:'ol<�f��st�j,��lR�3�0M�s�.�r.�c�r�'h�X��>� �b�ݦ#�p����N�L;Þ��1��c*eO*[ܫ�̓6�}��|FO�+�o^c
��x��d՗���)�w.�䧧�XCuRͻd�2dF�
�iJ�B_�R�cģUc�o���Q���䐳 */�ӹGH'���5s�#��K�)Ҿ��g��᦮9����F�o�����yPj�T}
xe�+�{J�c����=�I�
�4\p݃s��z�\��������,�