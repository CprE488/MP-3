XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���bJvi�C����M��Z�h-	q�%Ň�[G%�A��[��Σ�,R|���uP��g�8TxX�8�0�;�����Vn����=ӌ�{\���e�v��W���+9�]5.�w��W�#Ӧ�̋��r@��$w[�MyQFr�U��DЌh��"m�ukf��z"��8�,#�
,�k��V��)�á�w�P��,e)	1v�=�VZ<��(�٦|h`H���Ǯ�`��h�}U��Y,RܬE� R}6ylQ0�ٳ�� l�����lYj� -�ږ��*U"mr&@��.k�����e/E��E��I<VD��0Ռ,��8�mGK���?Pw��j�0�e�5n������)1��W��)s
g���x� ��`(�?��G��S��z��&�M$��XOC�ژ"1��^�cX�T�$�W���7�4���S0k3~���h�Q �!M�N�-���:I�T���=����\R,�G,�{��/��P��ıIh��V��E����=(��@Z��M������0h?�-�����|5aJ��H���}�9(��9�Ek�dS[�&���ZHR���� �)}��6�ü!lP�.f3�4l��.i�\3ܕP�q�P�Q��O��ɮz7<>����ٍ|�?hV���$u�����Qċ��=�v� Ǌ�ߎ��9;F���g����y��]�ׇ�iu8v��oz�&�R�07l���h���g�|�Y�����:���'`���乧�諴;��Z��v6�XlxVHYEB    1e3a     a20$�2z���1ԑ�XozG_�r��;$r7\�L����(�Oq���e۸4F����EW��0�|�@*����j]�UQ��yㆋE>#�c�4rdگ)����5���ϓ��6� ��5e88H���@K0���}د�%m<W��ut,nt~�FJ2����KVKC4���X�z���Mt��R����a��*�&fM�-�6�UK��ld,��֘�C!�1<�N5F2=�}�������Ϗ�`�� ����t�u��N��̙��	���p���[Xj����Y�� J�!3�n]��2�<���+_U0TZ����l��0��o�8�T-$�q��a�7��u&� lM喣���C&��lQ��Vg�T �Bh��CK����@�[�<G`���E3��ޏ�]�r\O���B��\.��S�����W�i �p����)B,bK�eٸ%��M����w}J?��������9nP8HW��6Mm�������Bэٟ��N�ฦfUʼp�0e�������u?x��s��Ԕ�Eud�(4�+d��6�Y�rؽ� �&�]2��\��@�*��9?5[o�I�E��ڣ�x�2j�h1?��'m��ђ�({���ܓ�Z��� ��S�!s�_r�j�+mx���`z����dH9!Ԍ��x��k�#ݲ���N�W���@�)_���2�*vX[��@I��B���D�����%)FA�4�Zʛ:MCfF��u!�*M|��{��tw<�wNn5����A=UӆC������53�w2�j��dD��?8@!�,5��E�m�N"s�l"�h�a��R� �K)1Na1T���!��&Q"Xo�N��I�@X� ��Ƣ�jg��uYG�4�r ��J
n] ϲ�t�qX�G��V����s��-(��~&e��T��s�kU��9&��zf�Cǟ�>��u~5`w����,�#?�h(�ѵ]P)M�	����`D�G۰
�2�FD6���O�M���Ѐy��+�[]J�r�:�'y:.x�L��;m�n�8�o��,��M�o��4���ZWU��G*:�C9�zbk��n	��������ëB����ÌO�َ�����B�����Y�X2����O�s�?:�K��u��?���l�6�����ӓ͟�O��a��l��qв�z�+�=��
{��R�j�4@����hr)�Cp��z�%F}�7H�ͫ��l�q������3�WW�1�(>;9����ә����N�҄+Ԓ�7��0� �!8�Q8��f�[ܰ���A�)J���Ȓ��	�찍��%&����z:#u�K�h7� �Xu���+�%"M������H1Nic�XLЮ<�Q�F�ب:�^����j���&����U�݅j�=I����o$-�`l�f��	WUJ|���f,ROC@
}���q��¸���Νv�B�	 w/�y8?��O�8^�%^KT��i�U�yCq�C���>�����A�@w�ucĆñ
�\M]��͸�׀:�lȓ-_d8H:&�>�� �J̴��G��M��%��b{g�2Rdl��������4�T��a�GF?L,&�n�c�~�MO1�L�i��Z�O(�x�7+۰�ͽʈ��-��v���� p5�=~����1�a���������<����i��:���s��,����;܄�cB[�ۢ�^����i2���&w��`�b��R��7�da���~�#���������?�Օ�҉���r!��m�bG#&w�\��f}�߾���Z�����ltb�ڂ��X +�S9��1����9��w�5G1�~4��6��.A������nGI�Q�V�0��3��sX'���׆U5"5�U\�~'~���ż5�7��t2DN�#}�a�i�==��6!���Ń��\�^��6q�u��'ZwGV�=c�c�������C��%������*`q�a<��	M�|Q�6�Cg���/xy��Q`�o�dσ�/۳��ʢ�D'���(f�7fY�ZgH-�*ȉ+�*��+;qEJ���@PgB����JZ����!T~-� �jTOk�	�Dҗ7*�lI|`X���������uS����4��ŵ����[B+*L�Ph���~�˘�G$˙-��9k�\ii�Gu=�A&��	�9ݢݹ��$�Ic�ڙ:��� NZN�<GF�@��a [�;ظ���L>lRhva���1z2��r.���Rm^1]��7X:�sVF	OIt���n?�>��O�3�X�x��d/<x���b,?�G����R�GN,����=�⧾��yi��6�����"���D`���=�`��D2D};�B%��V��p��HJ24�i�ҝdP��!�I������0��]ZU����ֳ�rC7�6���+ؚg��_-wI�	�
���#���O�����jYtzJ�>o�c̓��m���]���Kѥ�y�j�	�3B�P�q�bW�ƫ�U34� 8c�%��u�x�VO=�4���D���H���V�d�q��ŵٌٍ�t�[Ul
�F%���mP�*�Ք�Gd�����