XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����n�:�;D9,09ƪpv�Y����͆�@`R�Rl�b܇4wBB���1�xh W��Yǀ�I����^�<$v�Ն˃=h���wݞ��MY2�^��i���Q"���)�������F��k6�����1��es�Ԛ�0�'[Pf{��؛Pn�E�*����b�ԛ6phI�w􄲑'u�+B����Ŭa��+d{�>��:�&�����L[��1=�3�r^�L�ͪY�l}������wbHu�C[����2�X����!�8�!�F���M{���3X�qXxcg �	"y�S.1�j���s��&���}�~ 
�ʯ;/)�{ô�2�M
>{?Ov���c��ˊE��%�����,����g��M�BzfZ��>b����[h��W�U�ν�4E�i����
��Dz5X���Ȇ|��e�5͍���5�b �Q�rf>��/�{0�G�
���	ɦ0��P3��K�DFb�+�߈��m���=� ���)-_;�'DRŁ*A����
؅�R�/8�o  Bf���7������ȠҾK�@L�͖�Z)��&!�i�a�$a�@�����<�A�}�,K$;�f̑�'�(8��\g�\�PbOȪ��z��|�m]˖�+������n¡s>*�N-�Hێ�0[u��A2Q �u�4��j ż�|e���0�(�T�x�A��mu��tW�,�m%������B�+B�C���c�G$�@�q�1\�%w*�A6f[�q�ʑ�?�.�Oz�oXlxVHYEB    3d1e     fa0k��-6+�׫DS(��ɻKWt�\V���$�^�oR{o3�G'���M0j�_��P_�jFn���.#�` �Q���2Tv)�A��l�n	<B��ݴu��-��
�#������ X%@*��D''�nI��[9��t^\�W���Z��"�y�?I�	�U�eX����vg��y �����"U����g��
�/ߩ�T�b���JY��i;�C�1��Ns��1[��RO�V�+J�������W��^³���t�����փ�o`��@�Ov0�S��_�{=[:�Mz����0�&2{Ld)�8����7�(I<ܣ���5��I��7�Rs"a�4�R�4L��M���p�2!]���5}[���~�]�>�b���X �1����&�K������V���/��Yŵ��L���@;�C����ϯ0�w��ȓ�0$V���[Y�oY)��b]���[kW3:+�~"�ftW.��7���'���M�����N�/�8K�&����4]m:�����禋��� �5�]��[�'�$��F$h���a��L��x�U��/�����3�2z��F~tS�`�E�/�n�ĉ�������Q���0<%���xV��kk��Z��=)�9,�:زEn�NC_(�2�
&n�O]MIǇ~f`�8a���{�;J������F\X.�H�gz8jLG�b��(Zg<2L���!����,�.�l�	��\;��[PB�\Qb�����H��{C����D����!wΤ��s�4Z w+����S\S�^+�v�K��]
β .�I\�*�����	��%(}v�>A���h�T�J���!�0(H��;?3v�bъ��Z{��Ӟ�y��I���Q�I��	��2	~�9�_]���B��i��F`n�A$���eY.�d�29�dJ^@�a����"���ݽ�ϰ��I��E�_�(�V�#�E�"eVDԢto��^�	���I��H)���w�c�Yx�8|�h�*�mV��d��%?(�����l��C�L1y:U�hCU\S�+�b5,�IgG�#upP�9��}���r�Ͻ��g���,h�h/o6jK+P���;�8β��q0��%qK�nT����ꨭ>M*LG��FOZ�c��˞��ki!՟��ߘ��K��&���e`�����>�&[
��p��=���Y�X�B��<s��
�4���^ ��"G	>%��^��U�`KQ\����R���g,�:�OS�P��,��N�cR9��01D�DV����뾙��P&���B��
l��� �o��6����npA���.�����qIʟ3��W^�aI�^b�oh�|�i6I�}��d9^zP"F�b18��=��Z<`����. ��Nu��	��l��5�`R���C�;6":���	$�(��1�'�^A�m~ţ�+��U{ß�yh��vt�r�͋4}=�[��9�գ0L��J&�`Dk�sj<R
|yqN���G5�-GR�^�4�ǌU��qH\��01�R�:�cd~�;�L,��_h��S�LU[��6X��Xl�1�/��њ/���.J��sz�*�?�lvӨ@a/�0	E�����kHh>[�[��'��'h,F�Ų6�U�����^5zr�bб�>�0���6��(��P��Y^�����3���i%Jl���Kix����um�q��8DI�
���v�1�=/S�mf�U`������Ҝ�M/0���sT�����u9������6A �ܝ8Z���\�5����1����%YC�I`���-{���d[}���U��(��a�;���} �|�Y��:/�PRq^�������)�%�mZ>�$z�"<`_&���w�(j�>NЗ���L�6��d��U#�O�g��~���tu�N$F�R�-;?��xM�,.�cs��@a���D��2����������ŷ�ۀ����̇t�Ȇe;gF2(y$�K@�b��-�O־��X��v�������n��������v�3����7Ɓ���s;A�E�H�H{ =�P��n�Q���
 ��u��v�� ���Q
1V8�{a�p�v�� 2	A��4eg�a&Q驵�y[�	)>�,�O΀��ه|�MlQM����Ϥ,��v��khs�v�<��&���#��4P�����&�;��B?��K{N�1�;^_�)�J�#�ţ墉zFBN2�P���D��v*�p�w��S�Q�F���s~[��.���oJ�w��\~��U �>gߣGF����{��k��S����,��ut�2#����x�oU��OE9��`�k��Jj�t6��_eZ��t!y��,�������~��_��� K�0�BF�k�ƱEJ|�{��A�e�j���]lG��V�4�8v��r]�%�����#O�,+>���*4{.�<
m�>�Ӑ�xIPHZ���f�\�.|G�� ���t��*,� mB��p��"�u#��Ϩ㠐ﬢ��#
�W�umR���Ǎ�r�\ҥA�2��E�y7,1	�g}�r�~b�&�qt����`�{t�х�5�&v����|h��P+��ם����A/_�?�ؙ)���yPc��]��z�����u,G��x����"�ߕ��S)xO\94ǯz�ԭ���YP/���H#��3.�0D dЕ��M&(�[�vɶ�d(T1l���/�3&|�ZH�8�&��
d��F]��3�[,8"�{MJ�]x�/QY�t�e
���o�=d�1�O;D�ߥ��	�+m�%�;X�Ŗ?�c����L�o��ZI4R�[�uԬ����g�]���l�1�,��=��d� �>�:?��@�m���+
^L�j�0�o0���|�DjQ�)�H��FV�E��Ȕ]9�Le7�W�cl �����z@����~��i'�.�xl�<
�Sj��W�?�j�e6��[���s��H��4�ҏ����G�n҈f��`/��N8���2�9��h����NN�!qC �m�G�~-���s��f�,9�s�8� 
R�1�wޒ^�9.����c����:�&�.�g6e[I���f�i�կ]p|y���i0/�]ޫ�S4X�$v����ٙ�OYd<��ġ?�q58�~����ih��b�I�_h5	�T�ꄓYHz�*�,�Τ4:U�	�h�B��1H����v�d�@A��6�G�b��Rn�\H��/��8k�s�"�=i�,��]N��$�f"�X��f�*��~��()�'�G|/:W�w����p�}}�h�*j�����C�y8H��LQm�d�c.I[q����.\�&�t ]�yЏ(~����ċ{�o��g�eL�-L�M���O��6"�=;|h���C*��̞�E��U���Ti�.EM�H0r�R���[�Yf�5Z�T���/�L
Z�-=�rF�;W�������������\.�	�-s;yC:�N��vJ�v��2Q|�7�YM��L��s_$K�x3]p��^te8	6��j���I,Υ
��Q���I��Ю�V`�w�b��*Ą68{��VN��4�;���1�jz�GD��)��pΜ���%��Y��qN���Q1uC$Q�8Џ�)�9f6��y��v�E��	���LiA�[!�+�с�ϸ��W.� x&�'��R���&<�=-�,�=6W��c/�[N���8���[�a5���: ����=�տ��ʙ=�Y�%gJ���~ӟ����Y����8p�qY�4�?'�$�Щ���+�L���^S�&�L�����G0��z!K�E�3@���d7s��1�u:�]���ܵb���C�+.Sv|���c}	(Y�9Q4yR桠-�lF�h��u򋞨RS�N���H���>v㣾g/��n�;�]b'ji�>�s��'��r����F�t��["7t��l��F�1{�p��A&]���'٠��=Ċj�f�,O>%�Ӝ����M(m�ߵ[=�F��ԓ| ���Z�*F���~�er�=7���x�