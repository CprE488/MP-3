XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����$��x�:��E���A؏��$َ��g��1O�ɑ�.
(͚\V؀,�DzFn ��u1�h��w2K�r����)� � _�����S��t�B�'�����
!�D������A`鳓rB��٘�~c��9�8����ɤʘ�E��1L���g�	u�*%��`FSEd1)��Y+ID!x8j��������a[�oA�w릳W� =i� ����Z��+��V�籺�|
c{��^@=a�n«�-ԟY7r�:��+�i!�9��_�A������v�|��#K;C�
	zǼ%w�U�Uh��_�5�����W?b��0&bt3���4ܷඞ���Ǳy���Y�m�X%��	��/X6=`�0q\��}�EOVw�f�5��v�3_.r��t�J������]�F���\[�1?��3���ɗ���?��GL/�a�C��B��#��aûv��w @��G����YvY4ӞTD���L��T�=�R�.�Q^w�f���1F�F�r �vy@�u�Ƕɭ"��`�P-��!2@��aY���An�Y�ssk��,��#���� ��k(9qǶ�7�g,���L������;��w�`{%�d}߼�+���g���ʊ�h��!��ft���O�ac�ojs�M[%FcZLTr���>��%��4Y�$��#,9�)�L�.�#�&�h$�X�@�>Z#_�s��R+�:t�����r×�Kϳ�ex�WN����z n>�'$�g	݆6XlxVHYEB    fa00    2a40��� L�Y���!�*r�Mꦄ�`*�q��'R\�k-�o	�F�o|�/���_`.J����`�3�pt��m��>�����"�ju���ݡ��ùKwau�C'��nB?�o�QSSx��[U�u��%0Q'�q���`ރ�Ж]3dS��+D�W��Usw].�9�澱�����#���ﲰ�f�܉!�<.M��n092nėNs��_�d����`;�5�>��6t��V��MCw=_��V[����	+�����F�]��;%�Qҫ2E�T����z��6�I��`��.ݳ60m�o��>���=���Ku|5#CEi�XR�y6C���y�)y=
3��	��d˚9WeT�u���wq����~��|��rbT�Y}4���ފcE����'@��9	`�q%�Dӛ�/�BWڼ�䐃�V�P���t(.q͚S���6q�R��VL�^Lv!;��n6�y|v��"w��A��M��{[�@(�i)5b�p���Ҵs ����x(�?#�*Yr�_@��V��k�ɍș-j�#�-�=�%�u��I�;�"�-,̃w�a̼�G�ˡ�˻��e�q=��j]�X|��`MsF���aptg����*�P�IUƦ���<�+��R���j��@g��|s�_#�(Ţ��ג﷧N���8�8ǳ��9�<���r��e� c�U��q&�bN��ɛ�3����Qz��C�۸�g~�f�Ä\Y������^*�s�g\0��j{�f)q-���?�zG��<_b��0��ѻ���i��\�����yM�{�{�)��T��"�y�,�aL9�����A�;i�Έ���~�T��^-�B���ݫ������+,N�ɘ�_
��i^�3lɪ�&���4�^�?U��H�o#2���1��ȇ�����Ҁ?X�P6;�MJ�S��rشB	������64!I��1�	�:��G��z,2Z�c��n��?�)�
<����5��i��8���*d�Bف�3Sd����t���$l� ����ª	�X��팫���t�e����p6�C�T����D���X��Qik:i��s��ϲ���ag �ػ�!ۡ�e-��9X�)�nD:�e��..��ߺw�8��妶 IJ���
)T�>Ⴂ�/����n��8�B���OQ�KP�y����DJ�ݿ�*�v��k����k�U������>K&���(x�� H�U����'�xI�w�ޚZr�)C���E]9c�,HZ�)c���.u?���� ���8���e���o��X�x�A��4#�N]�]��c���4R�H3z�Y�R�{�;c�{�М����IV��M&�f�+�
�~z�s��a�T�b��2y���V�O����fTP)Ud';�T��������e�*�B��%5&��Qټ�Bpe��'_����0��2Q�
�׌^yC��Ύ��>2�(�:C�!��erwMs:���Z��� B$p׼!凱/ ��?u2�p�0�8ˁ��̄2�RVq!�Ӛ�#��8 �����Bv���)���B�UhsI���o�I�O��2$X)�2S�F����g�w��R��*G6���Գ	/o���2�M�� 7��c֦G����M����&�th�iI�L�eɭM���ߪ#{�[��	r�n�Q��CB�Dxf�'�����w,:`H�~��ւ��b�ν� ~ln�М�2wp9F�G���[��"n2���'��C�u����hqB�䎔�7�{#�T���C�\�c�R0��(8oO���d�ܾ�o^v�̼��(R�??s���md�%?r��޷����Er<+�M���D���������+v�l7��Q[?ʚW��Y����_�'��y73�翲��J�������OJ��\�:�U�4	O�S�U�^J{�&����ck���	o-b�ԉk�e��B��=�v����cϗd��]E꪿��$�_�����87n���x�8Q�SwV�qu�DIx��X�ϑ�!���źn�H��L	�P{�<u�؃�4z�˅#S�Y�w6�z��dڔ.z���E�n-��*����q�zXy��������5��x�`E��m�ݬm�w-��۾��4�����6�Ɓ^��B����#���T.��#��H�&��b�؞���y����٫�B��͒C��e�L����kry��*��(w@�SxU�$��K���\QVe�;�e�7��C٠/mzGY�'���$��7Q��`+��tq�U�����&)�I��(}kK�4�D<'�*3��p��_�HPO���Jj.'؞Z<rGFޢ-@�mR[g�A�����l�8��vN����};�
�Ѥ���#�:���|!Mj����ɉ��*�r��|� <r�d.�,��Im��e`H��5���C���7�p��~���� ���-���e2�Iם}�N;���,�[���M�����Ln{���o ��'�6�v����)��vg)j�R£���#�6�l�
qL�X��2�Y���B].�U�4#������LL�U��;��<0x݄I~S��oCD܂���ħi*#*�l����sK�	EK�N�m�6�.�1�[P0� kq���X7�~LY~�2Ux��x%���%S1�$����e$=V���&
�����gGL����W>��=QC��*���iє'��Z��X��=�+	B�˫k�kYu[svO��=펰���JB:&0�Q��-p� ƽEm�WD�K �{ڤCښ������^�p���G�k1�}����!���3�sw��%A���V��'��fР�����G-����XJ���sMt�2X4��5V�+��$��/�^���8� ]��� ��Ô�`���uP��}4�x��|x9�~kq;h?�0VAF>���f�n/%�t(.�*�Z�չ���8TVVo���<��dWM�f��W�(�j���}[(e�5�����M��b��P-�c!�@��έU��Kbh����B{5K@/�5X��QwۊR��3�Z��)�ֿ�2s����VZ�ۊ[Ĭ2�������n�`�T��9�=�у_`�j)�i}���/)c���j4�I�W�64���H��Z�s��a$��M�pP�MJq*�������Z�
'���>B5��UU��k�X��Y�>����RN4 �Q���O��vBuހ�a@u5�@o�ME鴝=�Kg��"5�l,C����f�>���'���^�ė���k��qu�l01�E�Y)w�2�{�1�2��}|V�ݽU���J�`�{Z��Q>�d<P�Kʋ�WK���#��Ĭ�r,�ػ~-��i��C%kxm<���&�UQ^��&�X���)��V*�h=s�P-i��a��҃�����p�A�b^)����:�b�����sg�aoDn�Qz��.l���]~o����l���d7�j\�,����ǘ��6�i�=�D�A=�0+�q���%��R-�4c?��e���)�&��Ov�~	�K��g�>`v��.ܑ�����",	h$�-�6{�vk2����-B�ܹge�c�hlD�Yn�+����Br9ژ\��^tʭ�(�N��:b�*CWps��(�,�$%�[p $Jp���/�x/�`	r7	�	[bA*�SUH����h�z�a��	��6�\�k�Zd�AF.$<����DRz���J=BM�:>�����aG�����B=�����)���W����
Za�D�>�C���qP�[�Q��ϱ�g����ӷ����7��?�˸�GX1B$�3��rQ�T��D4�T!3�	�2`�O��&�N�
�������n���A�>��;E��'�+3�i�i�R��U��:�&� B1��x.�(@�iKX�>�Ob�Y���L,u����D�w�����~�nM4z�=�Zcn>ԥ�|U��j�:I_TW�p��<���Y�����4�e���f18Yۢ�j-؁t�����PH�T�� ��=�J�t��w.%<�/���j��$�-�̀Z�?�n�QWY��i���@ EOÃ�W��5���t�O�
;�#ȵ��~OÕ�ϗ��;it�ԍD�L�{
�ZI��/���ܷ�m�л�-��ūW	�fzez���U���&d�4��w�4�1�ΐ���ɿ�`R��i�-P����KcG��
B]�(ؘ���J1����ȋm~ƥ��@{�9֊M�n�5ɖ9�L��{L�;�A��s;�QV���&v#f���C�,k|��q�lqP	����U��F�����D���gp��y��ﱢik=ǁ|��p���4]Î���s��M�;������qC��7��`L��eQWr���؟r��L�5��t��~���9�~�5Z�k˖g/�G��x{�qU	K	�7����G�,dr��gS�P�n�m|c�a`~�+�e7� 9�s7�<��	]�|�=�i�ЏM����֢=g�[	�ZñB���
�!`ܻ�����邙"�w6���Ѽ����������ː�V� �V����Ma�K�h���HgM ��l��}m�8�!�kbY��ʝ~Y���]|N�
�����	�k�SH�KD���8Q�/Ձ�����Nb��ܛ.W�(ZU����7��ZHL= �0<��-�o�red䠜#>�R�3rP6��?���.���6䇉��+�����_KܻU�䈃޽���MWЂZ1D�\;6�L!�l���#P���Y���%���FF�A���=�N4ѥV��e��fs�,P��&��c3:%�=`WY���<I�*�K�F�z��K�K�c������S�
�7J�!�X�=ݛ���91p�t[27#Bc�?67�� �J:}Yu�|���)X�6�L�,��Aw<7���k�.��{
k�,1�DG*�7�>���:��Y�$�P���Zg�~g9��7��[�_5��`������
���-�C���ޭ��+R�@b�cc����U[������~L(�6�`��8Z�`�u��]*C׌��B�ܓ�:'���(�(��ɣ�0�oS��#pܦ��d}�ɘC�̋�֥��+��h��FUH��`��K�_�؎~U��p�s{%5D�h4װ�8X�+�K(��5�ODKY�{1OrIA�x��� ����T��r�7��S'$��Xżb==OJ�vˑ}xp�@#v�3a�w������+F�����7��v����?\��1INr/";�Tw\s�t���5{h�3 !Рd�����B��B��]i����Џq�����UM����WVb�#a��9=��?�b(�붎;��v�@ʞLb�:�? ��*�o'��7�Hgz�G���V&]Z���ͅ��l�AF+��:o	�� B�X�db���Mي!����ta����G�Rz�j����TH���W��}�oo�.z3��k��vpV�d��@F�J<x�D�����#����?��L�;jG>޶�ܻ���K��Gӗh��g����&��v�͹3	v�?��X��.��x|Q/4�@)ɃRcZ^Jc�z����]��3-�(����=%`�b�����r�z�(�^�>���_����x�(�Jv��5Y����pX�p���(C��wX�����di�uU�J���vt���waN��3D`���4����]�T�(�5'C�X�f:����r�̻:��Je4j�g��P-�~��(�bA�� �d���g:����cY��^�!�w���(c��S�������h��V51G�R@쯶G�a���tRR.���Oo�s{���J<���^mi�{y�1;ŷ�T��X�v�X `9-�<Vl҉�����BhS�1�v��P�I�����$��t�2�B������`��p��@����b�@�S�C�$Q�6�A>�����P������`AVU�SKmۼ��C/��f��5�3f(�_�I"W��+�,���?ZY?
�ce[n��J�Y��"��qMG����j���$\��|E���E#{��Dq���&.Mx��'�I�,��,�V�^C����m�U�U����#cfMp���G���6NU�A7t�!X,�2PB�#���H�T�*V>�O�H���U���,�X��v���^:@f0�R���55�k��u��ѝ�rGD-�Y\�!F�mc�.4ɟg���ଦ;����K�ԗ+�Әm	��L�vti���Q�@�˄��x��ApAy�ǔB[/�<��ؕbܯ-@�7�,�9�H��z���
���~��;x�bߡ�!�,�(�w���(4x��L[���]��[���P�����>�6�cf?�i��k�'��p� J�qC_����SK!�������p@�<]��5��6�VԻ+�b���7��C�#�L�fF�t�R��Q+2�jG��j.&N6��aP�����7���I4��\���z:�_���Pzh�� ̠Wŀ�i�������� ���yK�`�]�؄��R���S��T��ď�Z{���;�P,%7������c��Kx�K[O����P��J$!��ml��'q�U�y����(����
êM��w�IRj'��B�O<.�i@����o�'V�Փ�՗�.X�m;T2�ȏv2��G�m�4Q�ٖa#+�p�2����ʊ(,����ֽ)XC���T1g��:K����,7@�bj�8|�l�$���At��c%�_�	�Y��SI�&� ��L�_]-��e���d��+^W��G�gH���=���*x��ALW��	ٟGj����}	��Pob뫰����p;,�q\����P�{��A�P@�'z���p����F���#>i�̬��ž�}�����㋓:�\ ��y[�q���w��D���:#�bl�|>�N�P��������_��������+���qI��pP���L��5Bc��X!A�����>x�U��M�Ү��۪��Mr�]h�g�_=`��J	=���ɫO��?���o�qM�MV�cy�8��$�zG\�� ����<��w�+��&��	�~VT*��,c�'�_q��ժEj��zfU��y��<3��Z��y;)���h���l�V��*�c��%��e1޷�bJւn�a3U�7���G�J�c��_�Ó9.�n�.0K��ᩕ��M<�+}Y1࠿��r�õ5��2}�«O�q�
V�����ݔ���O��wqz@�{D���)4��� t���G(�E�Ōz�OlC1��Qς��r��O%^u5-��H��#-�rL��v> O-�=��Z�l���zŃB&k��.�?�;�$�2����K3wf�B͑�N|OW���B��ÿT�9�J)�;�b��6C���t�����z�]}<-~�m���)YH|{Dl����G���KtL�^{��_>�Fy1�ʥb����Ҍ� ���C_�)�W������iZ�p�p#m�װ��E6�2?/jX'���̔��&�-���F��t@h��H�m>�gxdl[{N��H�јn|���hf��N���dI����\��fJ9a楶R�_���T��n���g}]E�g��[�GR�eZ���8-U�'P/���}oI
�dY���Rț�.B�(=�����4������g*��{}7� ��'' ��&��굳�Y	�	v�h78���F93�	f�I��ŇL�vˠRU��l����<�Ե����ulK��"�Nl����7 u�ؠ�R�\��p1h6p�agI��ҙ9�DD�{1;��Jx���� G7�Į�4$�5������~�V���BTC̳]�K����vO�o�_��h��ؿ�������Ti��R$U/��Ǉ�8�ni�t��yO��a���@$��b�}E�S�j8�F0�<t�j"+.߾-�)�T��1_���9�\du�[G�^��մ�^I�k���,ӜU˪��0WN��Q-� {`o�ڄ/|D���)5P�$�4D_j1��t��ކ*)d�J�q����ߴ[c�t�2��M�f�ם�����Gc��3Z�M�����L����x�P8��$���;4M�.����At߷A���<G�&�ڴJ<��hbg"t��ˤGH�"-�1�P1X�Zwİ\)V��u:�S���irB�%��m�Yb�S�x1`�KI��c�������R��[[OVx��rrM��X�����X<`����c��<��n�aG�0�B��t�7�9��1a�����s��:\� Z�wZr���b��I�����n�ŭ��	,�)�����X�8��v��V^�p�Et� ���a�%�㓒��C�To�X	f�C�(em.�����K�cKao�t�fy��+��r7b��F4=$/�l�gu��* ���J���sv4�J�p�&R���k�i�{`;n��8#���+��3���z+ԅt�GFw���(�~�"RI%pg�_<-&=��%?���d�e�-Az��*�JיF���3,�q=22=9S���"��K����t���J>�T�v��ht�"�����&�V�9�lo�|tX�a�l���ޙ��g�A��J)�ef��%���A<� E�!��uAKw���CPIX��׽Wj�l��|�_M^��،}x���	??�,�
�?����9
M�L5���̻�V
/n�"���W�d��s��iw��s�G�XW:F��!|y����F����l���G�%%7����q	�Y��:%j�nn���ᚯUez����Vc^p���&j��o�{'a�"�'���J̵r��,�޲
t ��� �^����W��J���;�	|I˃Gp�dQ���Yd��g�"�����7�Ѯ��ke�DR�@��x'�Ug�X2���f�2N�Ƞ���I����4K���0�r�	^�f��y���⣖�v�#�<�H���DS����C�������Z�����7�h�Ή�(�]'�SKe�xEkF�3ui���H;,��N��[�D�GF��*<Ώ��׷���Tb�ѝ+ȣ��G1�⎪���"Z5К��h�r���)+z`XM���tԈ��
��q	�=Jf�0�J�l	���d���s-	���K?7���-̄8b(r�F�f��Q�D�SāK3J)|���I��E/�$�L����;�-J�]��.+��Hqk4��x��z��#�5�8e��L
�8,��&�σ�7�77ՠk٫�������B-F�Q����L���l��EljR�����P�faFlQĲ@���J*���3���������Ͽ�K^kԮR�m�� ��mAIA���8���H�c.�3���M��>���d����P
SE�5H�-�
)-W�*���cL/�r|I�Tף(�l��� W��X)	�?j�X�q0��>m5�����%~6���zH�"�p�;`�Z���C�ln�r-3�<X�-��d�˪�q�M/�O�����N;�cLg[��c�!�Y�ltx �f]*��0������vFS�[�~�@t�R�No��,�f��x�u\���k]Pl�Mg<6�:* ��t��ot�Xb̿��:rS����wmJj½P�S��{�C�8E����vc�K^w�؆Dz�j�|&����'n��*� �8R��AUl�Q���O1��!�>����\�p$�����٤��F���S`<�K([�3�(��������B����W�_�I2���mS�&Ba,�p?����u�rs�& ��R�ϳ�J��4���q���T�#�f8N�����/���"l���lh��7����v_[�=1V�1e"�z�3\]�	Pp�9�y8SR:����.�eS-��)K�-3�Ԝg)w����adzq4�bUp�ȱ�kY���V���8}P���a�A�����ʸ%Vv	e�����0�g�A
^��T��tQG��40N!�u(_�7P���PM��Z���Ua�Ȝ�p9�1h�U��kC�e1v�J:k�rz��a�Ѽ^��gu��D˄�P��3L�1~�,pj��Q���O�D�<h�z'�0���:�
Fv�#��W��t,^���`=�����?�/��H���Y�4_��W)��Β	OT`m�NA��^������v#���ÛZB���(����o%s�|g��K�(�$���C�ɢqpbA�f{��L��H�Xgˡ���:��4�q��e���ƴ�����t�g����Z�:ey�Խ�Z1�W�9���l���&�ɾ ��Rٸ����s���Ra�ms
�G���_�"�z�>��1H��
�e!�R��Z�!�T#�cw��V���ꀝ9c��ؾf˸�;bD�N�<Ч�b(�\��G�����^8T(д�ّ5
���BW:���\.#��ً�v��eE�9NxI�B�����M�~y�SV8>���L�T�ͮ���H�	*���)���!��$�K�{�J4D�l�@��'NM�X��@�R99�5J*�Y�1�˭<
�nHVyޓ�"��n�B
^ʈ��W"L@�_��������ͪ�'�����+�̨�SC�5�ebV��H ̳��j����	}v73��q�9(%�x>[w#�N].Wm�����PN*��������5��/�����~��+�S<A�O�61cҿ�Sڲ��]��_wa�	��<E�DXlxVHYEB    fa00     8e0��'�-��b�[F���`���u�-sF���v{ͳ%qq�!GR��*vk��$�Cnԛ����q��D# ��	s���N�)�;L�q�.Qs�vMPK6�A�/W�ᠢT�SB5R�:���#��0����������

\Fs��yn��=߹�֣�}�[�ث�dʆ=��S��r�\���]��.O�|�1K��u��^ws��~!�ƥ��:�a��P���L.Z�-A��͝v�a��h�˂�۟��̳r�³��O��?�,�D4'-���[�ȓ�5̕�X���U>X�:'v����`W�ғ����~y)��c+��oL��ʅ��V�!�x�,��Z<_��e��j�Z��ש\�@Q�z��-q����G�٠Qv�g��`s�Ƒ�쿸s0�S�2%?)��wjꥐs�r�*��kQ�_�a��y+��υ ������O7����2�^ꂤ�9"��Q��G}aٹ��R�z�6�jbw�<���B��0��O��D��J�s�#��l�t�U6���g�����>�> ��p��[g}��`��J]K; �����?�Sq�?O��X!�d�;�,��~�n.2�C�3��v�!.+�b?��E��W��f�H�6��o ��u2�S�����Ջ�y!9�󟚀�=:!9���ru@���,��Vװ7����S0d8U��fٱl���Sἣ��p���g��!�i�' �-���F��V�,<���I\�ks�/Q��'R_�ړ�} ���VO��|	�ڹ0l�7*9�x�[��ߝ��OW��`m��\�䗷48�8����Q&"wQ5%���Q��5�;��}>~p�M����I�cd/�n�ؓ��nbO����1�|��t���J�Ϋ���{��ʲ����pi���ƴ|xL�|��US<W\��LE�C��E��j�8�D��>��O���ƀ���y��Jj�7(hQ;��eck��)��������{5ͦn�Q�*�C���x���-㋋�v�l���:d�8��j,�fůYx�;������f��$��=3���F$�߁@_��%��籠a�#�*x���>��wJv٨��z���6K�����B}�@���CT�h!���EJQ�Hj~�Y�1���l���s��G;���ވ��KX�Ts�.�j� ��h$�ñ����0��Sb��0um(�����p&�������eb�w<�U�����$� �E��륟	�)	������b��Ur��[7��xN�IS�*�g|_��i����>u����T'
#"Tc�L���'�a� �uCvQ��4��1����F�6����[4�W�|"��(Z����*�G��f<������s�}���㙿P� �h�[�Ɋ��e�@LiO�٩��/�b�zuG%׷x�+ҌG��S�ML��Oo:�R
?���A�gm*��1����v�TyC�"�#u�9|��������tH��[^�k�3Di����1���)��p*q��A�oj��%F��̹t��<g�|�F/�Z����?�� 4x/n�E;�z���	X�Ԅ�}�U�(}Q���In���I>U@%\�yFds5�����G��hTd?�Sk썭�ueJK��8
�l�����������1Q�8i]Y@�_��#gl��I�}Ǿ����e��c��~`�1�:5ݯ��廉�+IN$
F��t�1�@fΌ�*��<�����C*g
��˭�nA���:kb���埞K�M�6��r�y7�
;�Q�٨;�g6���Bdce?��W3�Ӧ=�)�Y�־�r�Iw�{5��*���]�7	�G�ܪ^#wU��ʱ�/D����q������K.���c���<��I�y�3y�
)��Vi4�t�թ����T��!��7zM��,�p�\��#H�!ւV��|�\3�Vf�G���F��-	3�����4¸�D�G���m�𫦮�>��j��_;R�T{_��Hr�訒�a"_A�+@�B�������NT�9��L�Z�?�"=�j�q-����U�K?��i
ԋ��B��B�?��B���i>���H�.��ӌQd;E���a��)W0֧^"kn(t�"5������V��������K��yh����}���c ��݋R] [+A=�ף�|Ek���|uF;$"4�| ��g�{�����a�d߱$�.O��M\.}��h�E~��A�����!<�tɃ�ѳ���R�&�_!%ϧBKXlxVHYEB    fa00    1110�@�H&���} ��|].n�I�����B I)5eɪ:T�p���S�`�=��1�;'��F�%�$*�ґ'Fx�n��uZ��Z�Zځ�{���ß\�ʆY��A^j'�[�'�+#�#����^9-���ϭW��P�W}Z�P<�ܲ��ϥ����ܒ����D��"��==\�L
!���� ��J�qn�By�%m����.
��[�^R����W&���zY"�r�A�-5�s���Gc�����H7���-�;�;�!TWo}O05E+D ��o���uj)�l�b����Rd���$�cC��pT�����^�rOf�~5{A��@s�T�= u6�c���(���v2�"an�/9��s�CTaUA�,>��c�]mR�������M��]*jzJQ�ۙ;�?{�&#Fq�:7G�������hJX~�I�=�����7/��a��/\J|
ޒ��-n�\�֣(�ؼI��oZ�~q���,� �\���p�  ������k ܫ#˄K�3i�`h�`ݼ���#O�Ԑ��hTT�BaB�w���:=�Vh���1�Ӥ+�d�c���kI����'�1��HYiߐ���¶��\�a=��B���9C�����X�Ԭ���r=3D=���L�������*oJ�K��z�D��9_mĮ��En�o4Ni�8�y� ��5�"�N��_v<����U��-`�4����tO���M����k�Z���t�q�a��|�N�9"�u_�f��ٹ��a�������w��PO�Լ�O�B�>�b�N2�"���ا��O�Д�X!�7�::����cǪ�]`�W���-�7QO��JlN{?sC뜎L�����c����g����O0����(�1Y��Jԝ���*�.!Ӧ�7��Ch�7�w�G�G��}A4�'���r����{N��N@b� �9�2�`VWS��w�1���A��r0��.__��wt�uf��i��$*6Ұχ���֯�v%�A�0�h>Ε,�[.zE��M9@!�sށ2ޮgG(��c�������I��|�sT+GѮy�-q�|�NZ��q��[�L�%5��0�^
ߦ�7L��J;O�H��l�'EBy�b����$��"b�G6H�����7K��r���*�/u�O�bǩl�²���Rw(��Mc��u��X�����n����D4kd�w���x�&�>�%�wܐ~$�[9q��?�؇�B?k��
cZAf����>��\����-�����l��@��r��I1�/��	W���ߕ/7̄�+�m�Rz�*/�Ҿ�R�us���!��,Z�F��K#� ���nvZ���Gx���i�E#E[%�d��x�D��N��U(҉�vym�`l���%��p]�׊B��7�=K�ߎ�.ԁl�A�}��_�r{% QN@Q
Mf�v��=�{J��i�Ka���H�d�{����倧��	�Z9.�Bx�jAܪ��2)���5G��T�*QԹ�O�Ad�'G���=h�")<�+FjK��ds�cOL�1)nvOh֤åu)�O��cghF��lÀ�f��)½�B���	�z����d��O�Y���S_;��Jh$���5��+z?�<� ��k�g�(��Pu��!�p~�^�2f�<��1�?��x�g�a͕�ᣢ��4�X�{A2���%�B���-.qʄLHJ@��O�!|����`#�rdRn]r3�G�m9�3�P]�M�F;髪�>�S�LK�i� +����L'��){:�L
e\�� 7*�K�c<�A;@�`��ϋ����_�SwP#]�ɵ��%2��ߔ�i{����9H��=S���.	?�%�'�;9��A�G�y���s�?��++���]7VOu����$P+���d���mz���1��] kI��d���A�xz�SrF'r��0r.pl���h�+��|l�&}Ԅ�r�c �ϰ���%�B��@��E/	�d�cY8��b�y0 ��y�$��G�`򜥵����5�T�~{O���K.���NP���O����|�Yҥ�y,�u����Y?��	�����L���(�lRgH1��fp�� �M��ޑ�,�͞~�@i��w�ۢ�׍�(L̖9��8Q��{n 'A|おE;8���H"��I~Rc�#��O.��J�b(�_�sA��|N}��s�ho��o��j�^c]c��`8k��a��:ڒ��F��fK\����MPH4/�&��j� ������n���Ӛ:a'�I,���y?�[��S�r`]�#_�d���d�p��Q�B�BVΆ�W<i#L>��^�$b�����J[��i�IF�A3V�	l�n-;�2u}!+&����yrV�U+3c�>�lK���|��D�gP���C��ͫ�u#�g�$�={��v������X�q�<��}��ы�?eX����~ *��ò���VU�?��Z4J8\ˊCB���.���D=��h�K}��1�t����̞�O���<�S���b�����u��Dl �1���;�&Vs�2�]�'��WE�f5�ݞ3��Iᴋ������4X���PG	~j!R���4�<4���BӉ��) w\� X�^��cA����ȵ��<�8z�!�����*�U�-� 7��CYO���>ܳL�yh���Z�C��w��@�����9�����)|}�l�Hd���["�|�IK����s M"�\S��x[{& /�?�ԋ8�ZF��X�f]R:�H�!^�[�X�b��B8��"&�H�)�ϧ�Yh��oY�M63MdL[�-���B���(�w��/�7Fc��p
 �ۀ�o:�1�$�^M�O�o(��:�� {ge;���g �k�.f-E����)]�Ks�;�?r���z��@�tz�Ci+����������Y�T=��{w�P�o������;�XM�g�D���9Q-?�E�^\N���J��<���_eE��^�� ���(���C�A'����n S��f)w+$qm���������6�A|�4��q���������|�c8<��R.�D�p�a�?������H�H�LOގ4�k�a�Ԇ�f��c*˩X:���LR��f��l�,p35�i}���w��V�hey���AǼ�pՔa��L��o3�U����.�+Qyz{�%��s��� ��DAc&�5"�tG!����;+�B(���l	�Kq3?��	��u�m�M�E:�����5�?$c��Y��|tNs�j��.4k�?!(M<K���6w�jB\����̻&�q~`�ycr G������-<��Sl ր}2�<�ǟ�b$��\鏎�G�Ԛ���><�ӞbB�`K�t�o!$�u�D��=̣f��&9��S�*�L�UT-�>-n��/�}'��?��(1�s��_TB7'����	�/��0�AL���t8�����!��ľN_��vck���K�r�5ر���+�h�bǘC����;�$��E��&y��ved�d�[��R�Z.�6��dr�vCtQ��Dj�G�2����XW�0�޿��맵Xa��o�S�:�1�;�c�1懿�L��J���oA멘��7GR�8XY$	�e�ۼn���(����k����1�^���M�c����Qk�Y	v�O��꺌��R
�bB��ퟔgfa��"�<�h�܃�$�;5+�����)�>�a]�:P�� �S=NI�M��Y��G����%C�aFf���a�YF♐����y�`گ�D���kPM�f��R���?D2�905kJdo�_Sd\VN��w�$w�H�95ʟ2����&{Bi������T�&��|�d41��6�3�QJw	�â�8�� ��o��L[z���e��Ш�d�D� �~~��˼�����Z����W�H����y��սw���%�q�O�'/۪��p�D�[A{y�{ 
l@��YE���.�ة���Y��0�wq�`�M&u�z@A��U�_f�Y�i���~�|�v��%�t��\�co�r0,��\vm��lSs�fz���F�Z�8���֭1��>l�h�Є�P�K���7��1K�KF�sQj�xGS*���❿���R~�8Y9z��}�������̶g
�ُ�<�1(K�zM3�k묦�����ԗ�1���U�ܧ�țe+�XY�Hi�(���MRv�+w)��m#��\U���u�f���;R*v3�L.��Ќ%�Ģ��iE�����CE4�P��	a����h�5���t60�{Q�o���D�C^8	/{�
�XlxVHYEB    fa00     ca0�ؓ���acV��8�*�,��lV���!3�	�O[1i(�=Ɋ*���@Ir�-��C9�fלh���e�)dC
pkQ�9_����J���L���pHz��y��ij�,>F�F�kэL�XR��񤌒�霼�@�3�ڲ�C6n�~�J|�H�r�6 o��z��s�R��4��%��&<j'�J�t��)��k�4*3'��1e9:����݂�X��Ab�<��h5Ux@W��%�WtΠ7�À�&��<i(�6�.��6��Tp�Y��L.��]�~b�ޑ��k�J&�)�6N����r8��Vt���|��?�!�#ا�2}��oSY�h�%������	Ƕ�f�
/���l��5�j!���옚.ˇzY��J;Uj_5�4�?<p��?{����I<��.p-dR]�y���[B������~������@�UU^�D�Ư��?��a}�u�)S����I��#�_��������<J{���:�|W�y�+��dg݇�Fs%��h!���E*P�f$�y^
�� X�и*����Hf�Xǚ���{ p'c{��+���`��
�}��cjxn-ck�cd�ò��z�x�
K��6�۲���<�Hni�-��!>�y�b��){��z�*/��Y�2��n!vK7�"��6Ć� �xqĠ4/OE#����E=/�}w�ӓ비y����g�蹺��ɻ��u�^��D�@f�����SmM���F`��ߪ�A,����58�s�'�S�vl�#6E��$�A��Q��ד�a{�_,Uou�Jm^�1�!�?����ӽu�A�B |EA��@����9(����`�9:*�]�/�eЩX����zG�O>���C��;1��O�A�f�pz<��JZ��T2*p״'�@d_I�������M���H���%x&ҝÕkCtZ����o~����ܢa+�s�d����-��6��P��9i���9v�郬���\W�7��[�P��MM@A���U��15��Z0�)�$;�Xu��v��s=�	M#��G�:�x':�������>(6Q���(V��k����S����b3 �-�3�W���a&��E�T9�."
�t�!֎�{\Pڧ�rq��(����o�H��2�z�}����C�x�R��3`�^�R��"���R���{a��qX��N������
��W��g��3�����vw��Jj^�`�\��-.X�l�.���8�% ���Ѳ�N�&"J�kiK�>8��J�PpIs���?�q���&ޡwEu���v�t� A�ϗWzOd��Z��TUJeK6���C���8�
�¯M�u�F�S�J�p�$����i���54��>]g��T�o]�&���u}m�c��yx\�Y����v���X�iq9�ǂ�3�� 	���jV�J��,����#z��� 3BU����@
����B���SS-.Z�GŐ�����	��w)/765,����Y��X�3B�B{vNr�|8��K��Q'�p��G��6�z��"���N�qkDs��\d�>K��0!8_�ifX� {�W�,sv9+ؒOd�|��P���0��!X����e�7U'��d?z��}��2>��>�����f܄G�2��U������o�����f���"��2���4�v����67/��AExi;�!�.#�EXt�t�"",ڱ��CjǼ߉�����w�o�"�w6h�h)IgI�2��e�y�� ���hs��2�f��c��J|���q�:�M����A8�ˮ�x��x�]B=F��z�v�#�|r���Y�	����
#�;W��\Y�x��j��r��:�ͫ�v(RX�%�u�����r^>�w��.�֎��<�YT�l�r)ߦls�W[M���yh2����J���2kx�1���@2R�|�	����A��TN�����A��_ކpٿ��M�O�Vˤ5�zL�ͪ�+���/B=���#>����M
�eF��f�f�2`K����<��a�,۪������f�N�s
�]�����%j�9_���̾1 V�!8��w���^���C
s�P%gP�x�0�%E����Ɣ&A�7l��sPŐ�"u����� F}Th�h�����g[@���3i���.���<ֱ3�n@\�#n ���,ֶ��9�-;�W�@xf�1�	6���'�����â�D��*)����S�6+�c\��HT�65���nAG���L�5Ӎ.�m�F*��i����(X�����ő���$�'(�����g��y��l�Y��¨A��{�_4�}�6	(v-��ֵ���,Bq|5m�}�H���h�(A�:Q��ɳ�|Am�q p��(�|�v�AYX���Ȱ� b����eQ�}��>�p+μY܎���E���mMQ�D�<^�Ru��PɏZ�ܵ[�l ��߭ۘ:��`�t����n`�'%��#IC �D���?0礍$�o_�O�|?���ܡQG�rt�1�ci���7�����W� ��%�i�͜Q/XP���¸���n�$��Иd�I�{M���V�O3	���G�R5?|�EΕƭ A��oM)��x>���οuax�TQ0����t��7oc_i�l�������j	J�&�_��IL�B��A�܏3��)�����:���R�O�\�K�����6�g|�Q�죇������%x塆�X �T`*�w��oO�#��)]8���UO�Sh����)�_5�jZQ�mVrEmj�����(5�=vHni/�ٷ~2�k;g�!��4�j�آHd*�K=�žR��\�(��M;�̠�y,�		����`�P� ���N��$oXm�'�Q�&!t��(�.~p������s��@�q`�9OƭGPHX5��F�
�˺Q�ݟ�	�T�e �E�!�s���J���bW{�t��H�fr��4�D��Y����?�d�c�dZт7;������<��׹����w��Mσ����J��E��Q� ���@¨"d���3�����(���Х#p��id����RA��%�I�S7
̈e8ȶU��WLQ+��H<��ם=�F8Lgb]�x�*.R_9��1�t��Z|�����i����1��m�Q2~ӭ�7�lA������ �q�:��@��kt�,�q�Q�����_��oo�@����o\U
U�~��XlxVHYEB    fa00     3f0����p8TB��ߏ���='J���Մ*�mp%��S�E���;��ՑT��V/K� �a����wS�m�5(&F�x��k�4̓9/s�q^��L���
�c�Q��Wo�Wf4h�hg�|�~�#x�������h��R0վ �o�^��F�AG�i6j����yf�I��ʾ	���rz>�-˂��Т)��I�o����thgoip�^_�aՐ����zC}/���Vf�V`Hڴ���9.�dX):e��X��:`kJ�����l["-{����8��g�3����D6,�N뒧���l�R��)��C,\�u� �Rs-R�Szh?c-�5$���nT��	m�o�t�e"i,Id�ْ�2#�	?�rSL��@�K�UF���y$�Z�||�h�4?��ڽ~����r})�(8��w�n#�f�C�V���r�!�1/�`�jY��Z:"�s��hΉ ���P��R���_�3���0��m)5�g&�����ûp����x9��d��A��Ex�)��T�f`p�D�[��hKC�~�>��ӱ�Ar.���8��� y/������U<I
�� $��F�#F$� �3�1���[U_RqJFs�� �n򬊽�y[J,(���?�����G-;����ܻ=��H�M�0PK}�s7��m��yIw��8�2����z��.�q�6��y!�a�E�}u1}�~m2�An���l�l�9�>T-YXX�� F��&�P�G+f�-(/z�e5��~�V����_�X0�)�=�Y9@@7��7�̥��6ܵ��G�2�ر��AM��y��7֛�OP U�>�n##�`^�K���vh� ���+��-R)lP�[�;���]���UK��n�ݛ���:�q'�%<=`�*ä�%̐O@���=.�0OD�P��q� !ơ�y��D^q�n:�����˘Ջ:�� 5!I�?�M�{��<Ol�M)EԦ�o�KhM
����`G�js}XlxVHYEB    8096     b20�e[^���o0T�����U�ش��MR�,Na��%�{��`�R�����ϫ�h�kc�N�S�J� @��G&(��j�$�ε/�1F�G4:,�i`���t���V��bG��w�a��P�Q*y�,&���[�E�������ρ`��"mF��bk��`�N��ǹ�_L<5�B�,	F�X���p�臘�r��%;u�3 ���{f7W�0V�AT��.�� {(��������$�L���规��216�AW��{�� #����8v֝ȥi�~�-|$4x��B�d+l���d@	�{��=��B����2�-�m��'W֊0!e���%��Eg��)���F�E`+���%����-�K�(��Z�� ��zTeW�((C��~�Q�0����E:`��7�`ogUu/C�L��O�Z�jO��T*�ا���h{����*ބ�1�d��e�*=����S�تR�m���3����Q5��KL�#>�R�33r�N}j���~��zR�\���y��Ԭ��������4�Md&���C�;�Q���r�L����r��I���3'F<c��u��q{��[B����5+0�06��� ���(,K{��~r~�k�|V�f;5T5�u
�_�|�"�x�����q��aGu*��=�"����0':Ѳ��j���q�0�v��$*�|&�����d|�����1�_b��B`#9c� ���j�����܃@f)X��X�x�~0�ʛ�ULUA�mJI�4W&Z���7��(�B�t�����j��V��#�m��87D'`7KIP����Kyꆅ,�x=<f[�����(�$f��=M��B|��P��~x��7�����շ��q�w�D��J�j�bq��!3I�4�v�zH�0"�f��`��"V��*|}m-'W�չ�ݩC��VHT�1\�2=H��ƚn���gW^A\R��52��׫xx�����~��F�G.~*NB�э��?�K'k��D��0!.����}�,gJ�la<�;'<��.,�f-I����cɅ�)pi�!�]���3�3G���<#44��!��q,bO��	ׂ�.�k��U�4�3��)��ӧ�|.-�ss�L��X�H֡$3얗���7b+�������/��]G���0�lY�!�^��ǿCg2�x�x�YR�������8H�ZT��g$��A��"���Ԓ!>�D�*0���dgo���t�M��砱��y0B�ր�'�x:�l�L�A��[������0ҧ�Ҿ�@�֊1b���c�D������f�nqB��bs�7U��#$�f��yh	�@v:�M�'�u���TƆ9�r�帘�HТ~�,h۹x0�1M���a�4BVTC׮zF|�����M�X?a 0op�|I�#9�k^�z���
��*��ꠉ��ު-�)�t�8��w��<[H�z�:���c0��۔���H��a�{w���W#�/�h\R��ۺ���#���o^�vY�lpt����]���w6�
���c>W��� d�|(������%/J9����`�$��ք�DB���Ѫm�8 o�]Y$MY�� �r-]\��F�����,��Irq��v �n+�l&�����ڌ�0�!����%A��ofd\�ݩr�H2�Wx�XG��k� �����c�g9��ǆ�ڒ�կ���k��Zt��`���\_,f��^�S)��f�Q�bW{�1f����"keei׺[�/	�V���4	`c���}@Ȍ�}8�O���2���P!�Lb��e�>8)Η���Y ,�un��V^((�s.��~Xv5Ķ�r���(? ��㝙[F�%e+壠S�r�X�k�	0�#�d-쐹C� +9Ӝ���
e����B�0�ѡ�'9*"Ε�ރ��Z�f�~��$�DCc�Lh�I�;Y��Ç�l�
u&�~Oի�y�l��h��;F�/�s��o5�Մ*/��t?�N���=�F�Y G�Z3u�ql"��5����z"���S�����Ɗ#�<V�ۆ�m�0�(oU�W��z(i��62jVN����B�����V�U�HI�-�t�׶L$���c�ι\f�*��_:�ӆ ��r]+�O,[`�����˶?겺�g��,z�e�I�將�<'�.�3�^�ȨZ�ݲ�hPJ��]<e���X5�e�����z�y���UJ`ܳ7h�a �;ʉ�mK�*0:��@
��$U�Dad��4�?��@.='��c 9�窸��-��\�Y-��E:�1�MZA,�9	[��i�"�ҭ�Y䵡�%����Fm�c��#<m�p��b_%����*����$AFF�^1�G��n$�Fb顩��i(5�����YKq��o�b��Z��)Z=�g�Ò?4g6|4y��5:���ԍ!����g��E6dt��!����o�L;�&$�iuG��sPzY�( �X�/����SO�r���F�Hm(f^p\��Ũ'�<$�L̑�N0�TX_]��!�d���l�ׂ �j�\���p�F���!u��<G@��9����h�~|O6Ą�,���*v��B�x��/���ߖj6�d��
w_����O�*��
���.�Ў/�1Ё2q���6�:���$���<�T{
D������N��f��[5�Hs{����=�����?���3�B6�5�FY�����pu���D�-��L^7��śt�0&�����L��-�����d*�����5PS�Pz��S��&��#�̻\��yYe��6�?\�-