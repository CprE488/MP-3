XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����]e��N����L�?�Hҁ���\'L�i�}�7�ƒiX,��"[]I�������%��&����!g���P�A�h��C���_�62R"M���ƻ�ҫm�������!�v��%�q���=��u͛~�ǰ�[��?�LJ��f���s}�]@G��n'��!m3Qzl����\��o�F���?����06��Scvg_B�P����"�Vڋ1
��!IT�V�Zb�bɫ.p`�Jja�I�����q8�p��M�d��^���R�EK^Y�R7i�X��b.>JA�E��b��(g5u�7��NKf^�o%l\h���.X�p����x�N�\.�ۢC=<��Q�n�c)�fҿx�G�x��\�;�l�v�e^�nsm(,���rC/CEǸ5 3��z�7!�^��d� �+L��w~��\�g�c챭��$��۷d^��ե����2=���Ld�oō�O�	�nxM���/����ޣh"�n���G&�BX���Z��*��D�b�����Y��C7nӌ�o8��d�[�6���Qꓟ��(Pa�� :9��~	 B�N�J�#u��h4+Sh�����	-u��^c�d�H���-�M#�j�����J"������Y_7s{N�<�F4������<�7]~�OXy2��<���u�}o�E�X�q���Z���C���Ɉ�Ԋ8	��q��va���a�,M���b �ȑq��p�aWuBy㬦�V)XlxVHYEB    1421     7a0L�lR���z��3��L�;��ثw˰�-�z�u4�$��l�V\��	��.����	V+NP�p�������$�)S�* �w(Tc��M�Iq�a~a��7J4n^'�_I5X4!��2�������;\\�6ړc �I@Wm������3ن�\z��
"2:La��:��hC; ���,��ˎ�<�aK#OU�ź�u� +��,�	�������q���.@g��
�n�sZ�T���H�R����DA�bC���D ���n
jte����D�R� ���gn�R��'!t$u'�]�; �^/����ןM�L׃�ɦ����s)n��)mP��K�)
{y�AJ<�n�Ly`МLJ8m���(������Q��C�����[�%��qw�#�})�I>��>m�&2s	�[�>��갴0G% ����b��>L��$�
��)�*Av��I�0lY�S��4;MzG��%E�)6Z�;N�B.@���C(!%�J�q���cz�ܞN��$ =���D�O�{�]�m��t�uj� Ӫ���h�{j˫��fT*PU�����]R�/^�H���p�����x�/R>���J��\�J Q���f��u{[am>>oV�g�yL���F��7�t�N�����o�O�"��0^'Y���D�x�^��ȟ�0�ws��"�s/a��,���A#�
���4�S8��#��y�Z�k�N��q��玍֢�Oe�ܭg��v��(!+2�4=�a��zE�b$��ʙ�9���)�=�϶�IN2౻ɋ&�(b���4�n������F�=��zp4c @�LN�u��IFK�F�7{*$�<�K���VL53�E�°�g<Sh��;N��X �<�V�(�嘷�+OL����~@cŀ�	�R��
)��Z�O��(rP91Ȃ#��݅��*���*j�Qf�i�@\]���W1k+������<�q�!w�,f�e�
Ul�௩��U���P̣;W����X���6��e�J�+�E��>9�؈ߐd .�� 4@��}����j���+7خ%�������5%�H��Fr�+�v����[��I�LV��n���m�*��{����uHH�����_CGk-���6�.���a%�� ������8j~Ҳ�N4G@��]<A[~]�V�F�.�&�VE�5�&C�vq��P�����!��S���;H�hf��(�ۿ<gWPCO�.8�����K�
����}:�� +O{�E�1�@����(�˕�F��,@DQCVA;D�_��M��/�ŌB�OͿ����~��I�`%�����v� (ii��&4�E�n�u+H}c�������Ð��E�=�b�ٔyz��|Й��I�V�~�J}�T�\�k�Y���z��7�NA�m��_�����-��+�`q]N`����~ ߖ׉v;&�h%a�������N(Q?4R��{�0�EE~���ҩ�`�&�V��^6��$�⊘b��͊�����ړ�/�5U[���Ak����-��tUХ�G��w��3�(\�IvG=R��iz�(�|&_��}_��g	r2\Ӛ�v^MS3酁1X��gٙ<�����"݄�[2������S(�k)[�i���!ݧ���רlT���A�ES8'��#�~����)��.���GX���\���ː�x��X��	����'�V��Ƕ��>E�y�hs6:!�Et\�W�О�Ϝ��:C%a�f��H�
@qhmP:�&���$�p���;��sp9�/����P�w�y�r)G)nO&�]��AF��Y��F����h@�v�c�y�Ǻ[����OT��}Q�U�r�~�1p �fC�V��hn� G��܃�`L�"�O*_^��ݬ�m1h�\��6F@ߞ�#�=fg��8w>l	j�=[h