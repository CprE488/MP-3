XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���W�:���F$�,����ՒB�Ei�a�A0{3Y���cN������y@�$'�El�w��c2��Z_e�Ė��,�O��=/2H��Ke�P��Ɏ��ŭ+FZ��M2�_��� ���J��3��'���+n�lO��L|vk)��ӂu�t�U�g��K��Z�C����fR�0�{`L����G<�X�"i@ҢI?~]�ƶ*h��|u�,^�<×�{@�X�5��c��'XQ�7��!P��[d�����S�5��:.���1'1��&���-G��fm��m�[�#҅���lL�A�:���VܕyTvLIs��l��9|��$0��"� Vr)��i��Ox!|V��Fs4��(���)�]1����&���
D��Wk��͐Z�#��v��i����}�+��k���D|�Ez�-�@k8�����@m�DlA�8H"�E(%�c_8�O�kf)���GӼ�\zP����~�Zd�0�ф��_+A��uZ] ���'��C�Q|�S8��֧w*(�VQ���ֶ<3��I��"J�����Uv��gׅ�CëBF�3�"&�����Z$���������9dU)�J}�_axZ�pIe ں���YX��=^�4m8�-�0̵��w��mU	@��Ra���5��Kh(��P6�3���\�Z����O�Jm�F;�i�ݳ���m���>{��{�]U�ηC�3Q�ְ�-��� �8[/�o�~�ݝ&�@�aeo~�Dcټ�QBM��8�S�u!��;���XlxVHYEB    17b2     880n�1Ä`��[�Ulp�m�ǝc�����6�eh�\>��iy� ��q�)����=d ?�#�^�ۊJ���h� �ڗ���p�E�-i�g�zQ_ڹ:o�%պf�V�X�m��<Y9G��2�:�z}�S���vy�C8 �x	c4�)�=�.t��w�w*�L]�v�h�5i-u�u��>r�'E�*�"`6);�T��c.�kI^���-w�����Q���'�K1�n���F�y���R]�����d�I~= ���5me�.�<]��os�h�f5���8�^�i��;�����~Z���%�m�7
���T׊�l#P�C^@Dc,�">��pt+�]mC�ы?����~?����?�opQCL�<�}�k�}O�	o�{��ag2�'�n���������CJ�A�lWCR�%;�%�{ߟ��s�{ۡ�lTヸ�^vv�g!e4�3	Gyv�%m�\.Fw,�n2�`��zp��'�*[Є d����e��H��/���B(A(���ێ�m�&���(�+�����lz�!γ�o�lK:	NG{NT�䃯�X�<Os�3*$�W�v�m�����]���.
�Y�N��x�zU���Ց��Ь�J"i�|co�iŻ)-�k�!�O�E�*x_e��^��>2�O!���g]7{H���
(�=	 ���tA�l,��������7%��Ms	��Z*�F	~0ߕ_��l:#Tܖ�T�>��d�{��ؐ�m>:�����Tϩ�>G�3���x9e�|c�ue�^�=d���$�Pn�R���31��� ueK�#c6���>XH+����{��B�P�����x�V�?�2��Y�9B������ޱ�C(G(��GS�n�1��h{�n
b��ǹ�j`lX��C�r^Mm,��lWٻ��<!�BJ��W��:X5�/�
�zn)�9S������N[y�
Zi��>�˂�@j��0oM��y
�:z�(m���OSC�O6�0�_��5�loG1$��u�Mhs\�Z>Z�'����GY:kl�$zHϣL�:ڬ�������ϲ�Se��4Q�,/���p�P=�dz�_>H`ft��m��*�c���M���b��2Ý?��?Ou��:���B���r�8v]�3�	�=O;�S2Ѽ|+�O�^�KIi@U��6��5C;���F+x;1tf���픁WΈ?V�.?��N��B�ؼtՇV*]�I��V���,�V/�Z�T����S���фd����`�q�5/-��p�ZB��E�ɴ�����a?�g��W�B�zi��f8���
�B�ğɫq�eh�E�::A���r�����D�*���@- ��H�������BO;2TL�<ǯ��������1���y�)����+����k5>Ө���l��m���A*|�P���/���ЉZ~���Ҵ��>���Wq�J��؈�@f�y�oY'����A�o�*?cE>�c0��q����}z���j.��ʶ��&��&�SX�z�D�����)�+Z5��z�9B�H`��ҝL$�f��Q���y�OV�!v�1�YG+���Ή��"�)aWsByAP&�W��y��Vw���;i$�%�
^)��%@ύ��PӬ����"a��']�3aqI�k��9%��ʖ�h!�K��"�)�
�C��<�������
�F���'Cz^�x^�@�QA�5Ն�G��}.<��6ٜ�}�4\g����T�}���J]g@�P_��$H�A�b���Q�͔놈���	>�E��� ��:Xaߠ���]�Մ��1H4&��l~U>���P7�C���;&����o�gk@qc��E<�"�mK��^W`^����^��/��7��m����� �r��yD���nu�M�֞_E~�]n�ݚ`>|!긏Tr�Ac�<k�/�\ ��/L��"/���lxJ�}*?�f�r|�ֹA�W:�/K��`w���{��VMY [�L����F�=����XeuB	��w��P@Xפ(��������	�$���remřa/sw#0E5��<�m�!��]1�|��G_f!�/�L 4�;#�p�������q+�3G]$b��$�U��#�.�o�Un�,��ٺ%'�����8�g�W