XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'�@[��$���,.s��R���A�;��|�?�`}���KlE��(�o��l������w"��	
�6�0���(��5�y�n��O^��2�P����JY@���Ԗ�p���s7*W1v��u�"��V���(���0�a��9~���`Q�<�<G�Ȕ�4>#�<�9�gR��'��7[y[���dT�S�|&Ho9R���P��l&W�R뫗��������F�P�s)���3�_�@w��O�-��R!�'20��A�YEÌ�8' ,�������65���̒�V�t�|�JȔ��~E�w1/��O��ž�8JzR	p4>�1�e�?+�}���p�]�s_.M���A�H�G�&�U?MB`�a����̀����oʪv .ո���+�^$JtȎ�Z���a"�c\�����fV��u�h�|���@����N�|�0�2ս�n���`��sJO��BH���������Ѽ4˶C���v3�pyXr����f[�ڈ���/,"B�9�Ay��&�3� 2x��J����L�ී��k(YQ/1n5�zY\䪧Xo����	��^�aUk����;��	���n}�>��y�^�)t������1aF�#��ͮ�o��
H�^	�عBL[O���K�K�}1��,����7�������%��O��C�	�^|�$0��%�L�r�� NU?>m܃�42d�Us6� ]3���T
2�8jQ�_
���m��|�v��ȍ���o�V���or��.N �XlxVHYEB    241a     ad0��9)��$�ĜD���bc�{��<K �ωW��X��M�����/��q0�̞�uQ��&����2���&�i�^�����;�#�az6U�b�Iُ���J���Z.}A������߿q[6v1{�G��2Ol��gml��n�q1:�%rl��() R�p��5��F���f�bL�����8G �+[{�_`ae��|0WJ��.#���4`}?_��}�S���ؽ�X=�i')���B���B=������L�Ҝ� �~ּU`�#�qHk ���zgq����K�A+���m(��]�|�i��m/NR�}��9�����>ޓρ�Uv���([�����.]�Hy:6���Z�^��4�=�^��~��	*#��Fe7�[0�A+�0�eQ�5�҅����`C0�X.y�l�~��j��c���P�74�L��2�\�屏����L7�6�}���11���ʽD��#�E?4f�c��r)(]@����H*���/�۞�G�.J�U�O]KH�'��|0��R'�ٟ��3x�'���'���kE�L�P*�^vP�?���0�g�!֜�K��m7�;�F{�R�2K:(H��YL0ѡ9>� Xbʱ�j��e�R�G
�+}G�����,!:�(tV�Wuq`,�#Gz+�j���{�>�����[�m��D��+��a�g������w����
֨�����	�|�eӲ}��6��҃7�؆�����~���_�ki��7�C5�p���M�� ?�X&��?!�A��4��2�r��"�Ȱ%�<!�}0םH���JporFfAIB���>C[��ħB$<�� I)큞'�
�i�L��5[�jȦVwD�L���Qv�A&p J�Q�� ���LB�{Ԟ��ǰ.f~�w;rCT}� ���hG�<�|y�ʀ�����Z��'�3	*��;=�����:�5����ʵ?��e@v���� �%�֢�#n��,%���_�V@��p�	R4�F�3	����][X��o�Z�)�6{��$s���:l\�$�Ehw~Tv��M,k�n�ģ�n{�X�h���I�K/"J�=d>-Y �|�lO��3z�KMgz|�g"�������w�	�O��eG�m<�~u+��qJ�-#��\�'�����\>�u�<��ˆ�tQ�X��Gx�k��~���"��9.N%x�{S7O������V������1}�c�,p�۷J>,���y���Wl6�y>������͸��)v����c�(µ%�!3c��e�ݿ�uGJ���uX?Ez�̰�6�� ���8���G���;$'ul�wA3~�|�L �~�'q�,nqr�:�X��y�r�OtE��'�H��6Tq6/������&[�#E�؉�
<R�t���T;l����s!�b����K��	@���c���K��ɭ[���B��L�=.DQ�I{��G�́��5�}�r���\�`ot��8�2�=�O�z�	�9��D6�
����_�EV���<����zKf��V�e�~�bS3�4β�6�Ϸi)��г��*N=�&C)�E���#��b#�V��ȳ��#=2��Ţt��G%�̫��Q���3�����(����I�����\e�sW`F��	t�ۈ�."<���`�j������`÷�s���
�7gd���^^8HN�KU����n�%�rS�W�'g�a������aZŏ��� ݵv����4,�hˉh�Bt��Ԭk"�"Lŋ����H��+״��d;���xS�=�ůʩ�(ݘsns-xFҎ���nd>�KJ�������=x,�!���#�}�,�'�U��&A=f>��R���V��ۃ7`K2'=y�{V�����H�D��5�'���C�����U�Є
�� �լ�{�P�����x��e�_�;m6�i�	�~��J1�CxG���8\C�Y�Zs'��g�i;�����I��2s��?��8�x�*���tiF�aϐK{	���Gk���':�{H~2s�㇅}�<��Ua����7���9�/�&��u,�T�'�`�`���Ƽ�Y_���@W7��4s�Ym31i�~W�⠗�A?��|�e�%�:���E�6VC�"�R������/b�]��d>e�GA�U'5+	�Ǻ��ԗ�h	 �5�D�#;�7�L��H���k�U�Hx�ҝ��c����-ޔ�n����WPk58#V�,ǣ&还���;y�����>l����UUa�<�2��Ý��Nb������cK.p)+����O?�S���d%�5<T)��f/��FK�mq��*�`ݬ���
�MꀟB|w��<��%�֚b�V͋�8���[TBF��;u�4ƴ� ڦKL�/�ںp|]�&غ����P�Q{����͹�sJ6rR�B���Y9X�o0E]��=C9�U!����
�w�of`�`L��0vD�u�	+�۪�٬s�/����<s�O>�V�U���{oӀuUG=���Ԇns�MSP��LW��ռ�`4kF3��0�1(�F���$L��f�ܷ��Dr����{�W�����+��ʇ�����G��c��(X��C��CG/0��%���9I6Uz�����ǯ1����6y6��lav���+n~�F/�4ʏ��O�M٤�3��P����#� ~�bN�Ցէı��|��Q?�O�7ƞGS{����=eK(ŝq-�/�A�߁��