XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���t�>���k]-A;���@�ְ�2�/�������m���w���-/��!	f�8Bcx6��1��96�?��#�4�KtR�nH�'�/F�NqT�x�M�n��%�_���J��dc�Յ�"N&KL���	���N<h�Zӫ��C9��ӄ���;D&���\�ɼP�.v�o;������xn��2'�x��2 E�;������"��JP�d3����f��#�����$w@���j�9�k�;M���=0�L�-�?RG6ڂ�3��,�
���|(��|6��னE\fC��WūE�´�Pë��!-�gr����nˠ�x��B�ڭo��D@*V5���xA5���\��s��.�s6|�C�{���5��:�-%;�����wJ�.s�]���W���,�l���X)J���)0���Au��R ��k���zo<��d�,��&��'V���ҲRS�.\��[%���m	������Y�u:^��	T�_q�����a�E-�~䝳jc)���r�p��h�&2��/�[�L�Y���6�l��O�e]�In�X+M�'���gj)8�q�;�V�c��h�C�.��{�k^�V�ˍ�w�i�����^�q�G҇كt~���U�g����=�����Z����1ʠi<�ʞe"7R�;�z����,�!���":S}��[=ZM_0�^w#TT��O��2�� �,Q�,U�l����A�8rh��vx�gy�,[�瘪�L@����"XlxVHYEB    39de    1170��.����H_7f�s©t��x�(���j0ӡdX��E�g���Jy%t�nW����ݪ�z�B�[ןB�o1���=����C�|���~�N�I����Wl�����u��k�|HN��*&�k&VF�/�顖��ޏ������fjb�R�}n��K�x��D��K���'�8�)�-��&���),�����S��=xۛ�h���-9CWݺ Ś��׍$���h�!������*@I�Dk�o{�������i����(7��#�-��׻8�p~�S�����W�5#���>�2���\�O���+�RUs4����#���gI��	c��r4�U8�7?K�\��Wf^FU���)��f[�w
A`������QB����P����� ���2Y��Յ�#se��\�@�E��NY�S����*�W�H���WPe��8/���Ϻt���7��.��<� ����WC��a%��ѢG��fK j<aOj�>��!ZԷ�>��q�=PJZM�O�F�m)�s+x��.������z�����o�c6�����T��=��)�P��
��e�t��'f���[�������v�����NX�����ݥ9������7�w^��O빁�t�,�*��'�7�GA���U�s2#�/��|���fm
�z����Pw��a8m�q1}��
����l�*?��?q!-����QvT�Ϊ��	u�*�9u��u����o�ָ7!��5"��)�M�Pᶑ�aw�ק^�[��K��pd�/�"�F�c3B@�R雫��'.��a��/�Ky�7�M�N3��i��/d"���Z��ɝD��Շ��A^�`�a�O��(>r��K��D�5�nhԊ�V��v�[h�!y&\�;��b7�0�"�%�f�C"�QاO���b�� Y�s�{�!�7V��v(S�D]��X��u��a�~�F��{��n�OT^G&����%�f�4����P��������aSeO�o��V`ʔ�!���4A�W�v%Q��Ȉ�C��hw�^R+�րV�r(���ʙɢ�=IL�h��Ň� �f Cj
��:�S����f䐄ls�y~o��F�#� F�� ��(�� ���/��u�5[������A';�o��C�(����V�Ja���lԹ���-*��B�5eqp5N�-A�1HW�\�&�cI�.w;����$�x+4�,�N���g���=���'�z�y����4X�J��S�Ղ}jnN�$�_�Yl<���6!���7�5� A��US*'/��a�U;T�ʻ��,}�K��zZ��5��z�D"�fG0V	�[�3��L�_&�1=nQ9谣u�ϧl<y�h��=a�0���w?���(��i���8q�&X����s��0��'�Ӂ
YY����nt!�y<���r9�cѮ���7핓��F�sq����_�E�{�8k�\Y`~�7��R�
�MO��`�쟩��$�}��Eh�ȶ|������-��)
����W���8񨨘hV5��yX�|�>��Cp��&˾��A<�	�ܻ�F�Yo��)������rq,T����~S<�`u_���W�V]m�-t��͖>[EH�GP� b��Mu"c��哯�/���I���֛n��]+�
ߧG�.`���hkʎ��%%,�o}�E7PR	�PE��`�;3sS�C3�y�I&�b��iѰ5bu��	A�h)Q��pdu0ơP"�뢌&<��g6��n̠�,�k�o��P?���=��B�%�An�%����hgڮƱo��29Y�m�D���~���qQ� Va�8�bb�n�C���t��ugkX��#�`�)2D����m!SM�T�-��&����xs��R�M�d�$��/ݎ�+��z�T g3>��tH'�����@+p�"�_�Ŷ:2��/�U���Ȑx��T��Xd�O�S/p���\��*��M6�ڱ�$Һa�Y�S5�aEn��:Ҍ��̀awԡ�1j�]I�Kc�?�0X<Ǘ���'�_��F\��:0�iV(��|�-�m�3��%р���,X���]��v0����o:g����j���`���K��>��za�<�����!�T�����um*ڡ1ੱ'dV��'����/��m~��x����@)^��L��}VN�� �J��%1�5���_zʂ=��L��������	�
�g$� c	)OqF\��p�O~o�S+���FИ��R�g�7�8
A��L�������iA�P	�f�Ė=&��I�a�[�w��������Ò%L�"�ĥA�so{9� {\u6�D���;����iP�Jv����^�/����0�AC}�OU�SV<-�u�����>uNܐ�f3�FlKr������D����@�:=*�%�	V�	e5�yj�B2oƘ�j��ƴ��d��p�Q��b.N��V�3��⼇��� �	7�������n�л�D�loϝ�E	��P�_2�"�j7��N�,��כw�d?�e��ջv�È3���N�0��4b���^ހ&�ұP�H�3�'v�Sܻ*?��^P�dOE�=:u�L&Lڦ��F���h�3�C$�~����i<ӊ�d�ѕ��wB���+��e��E(�Yd��'W���b�řj	�����C��Y��MG+���p��4u\tQՊj�q��X��5��Ѳ��r՞,h�  6�o�v�6B�r�:�n���6�}* c���z� �<DMy����i1<ӓ���2B<�7
�W�r"��P��� ��2���9�|���������0H���F@
�����o%��aˢ|���A�h�&C2�ְ֖	<��7:����-���{�K�f�#�y����o"�K����x��?��|w{��Q�#���4�SL)��s��	�=��8�p�
k1�/[/\�Ի}�+��+/g*���������Z�1?�f���?Et�����?��!�t���>J����W�>�� �Ɓ.���ux��}	�}G*u�����b
��.��Ѭ��tz���׵���jv+!1Piʭ�T՛���R���r�R�WQY{�v��2S��Yp�����zj^6��zՍ���u"�H�D؍�� {�S��-J_�s��k�8�e2��^?��m��$�y�<���bd�a�z@x��'y^c:v&.�Э�$�lSPM�!+a���Չ.��wEű
c�����5�+E�D�R4���M�0����V��9�`Vu��gK��.��,�xY���Y#��>[K�N��W�hJ�(P� ��n3ݶ�p���`��~�"*/��>N#=��e���PE�!����Jl�/45�dDw��1Qe��$"b_\��|���׭��(�8�б	��T�����N��pO�;`��o�z
f~��/�e3k�uǒk1A�|����Y,�0ڿ0�@ԫf�u܍+��>�}cq��J�H� �GH�i�ŧA���	�B�쑊؝�"���k�DU5)���I��Jh�e<Ę��i�
�0T8��Z�#Hx0�2u�'Od%�u�l�YfCjfZ�;g�R=�[���#���Z�K[���qu�K���[-L���ќ7�v�=�����q �i��a�D?��T���d �<�8!FHT�#5��(�NΔ[D�Gٷ�'�:<�z�ml�O6	+�2��mBG;�Y�/B=���Y�R0Ժ!4zA�-]��m�� j|l��T�#����Z/ԂV:���w�|�O֥�k�K���s�{�r�_���]|����5E��4�ܑ�p�6LN')�$�O�}Ä́���=dG�����Y7�ZW�"�fɛ��l��W��*'��L���po��ڒ��J5i�EN㞂Y5�w�q��V:bq�ğGa�@Y����Q�{AB�aˈ�{��12�d��Y�jw^��B+��'���-k����~o�>� ?��Y��:�׵~��3�}�ݿ�u�JT�������ΰ(n#+4��H���y��ha�:rCsD1-Nk����/�)5~C+x<��ˊHDY�q
�`'���i�sQ�We��=��=%��
y�xj��'�æ�y�=������[�cjwJ��wXk�v�`C� �P��+�z�H;�rJ��n;NR�-����B(�.o����NC�Cm7M`��!N�-���˲�Pݱ�z�O�c�_|LO�a���:�bC��E�eG*�Շ����>�� %�b��
���փ�uGGG�7b����Ǘ�`���C����(U�8���._�:�1��x�.��i`�� '�M�_k=	�e��&��8f�UgC7�Ti����z��I�,�;c��9t.nHb��M�t��4"�|�j��_�nʹ����L�s�Q�`1=\:jOT����G2��3,
�O�2'�&�}(