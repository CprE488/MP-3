XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����xܯƴ��|,�FV6�ƍ�fO�q�
�HK������ђ;5<9��WZ�]�%���
xN�FݐW>?�ߣ�,�[m���
[�&�]��k[Va�=K�K��@n�R�Ny���aR~�0�^/� ��3�Έ���n�>�Xa!I����Ѱ�z	+S�6�,����y��>T�;���JW�8K0k/`',4^_�Ҹ��)�0�P4 �N�`��BAvI(nQ}��	GȃްӪ���X�.!��|�D&�Y`[�dݸY�m��p�kFw3l�1�r����}����ޘ���A	��^c�Z�Nqv��#o
��m���J�%:�S��)��Ӻ��%���[� ?\?'�9`�u�D��7�6OW�1"Ͱ���� |�w�\;U;)��A�!�8y�j�5���=�W�����,*���E|3E���Y���5E�)�59ai�o��o쭍}��Ԙ\�7K�H�\_V��	~o�����dWAg������y8�Y�����D���rRO��sɊ��v�x�ɂ��|?Bݫ'2�x0H4��ԛN3��36Ft.Z���	��𨜝-�T�r���Ģ�Z'���
�Md��Q�}��ȟ����`ƇOD�p�J�3�� p�g��|X����f��8��L�	N��*��S�oE^0���^�T�~�J�y|��<�7}� )"�C^gJ5����]�q^Ĉ�+S4\�9�+�eu���ZKʴ����� RAZ�^�(vz�;:�J��4� H�4�1LXlxVHYEB    70a6     b90+u��%
�Wk�'�DJ�b_<4�����r�~r~9�sA��
.?��* �z��i�"a6�N��E0��)��I��&7���=q)���-��r򻉫l�Ǩ���� �/�8g�o�?-XI"�kMR�ZF:A�u�<t���*��]e�n�����2��ww��O�\
���P"������O���<�Ϡ��Zq�_�	����Ff�{��ĩ�����頇4&݀b�E l�a�#�����Q���N����Vw��1�9�N��.R�C�f&O$��ǎ�~��Ţ����ڦ�$��i	��p�å����]FV� �s�5t#(#i$�4	��t��t� Ϩ/B���j���&7�h���H�k�"��n�S��AR06�+͍�V���5��9���'*�?�e�N5i"�y	��Yh��e��`�5c�Nl�4�+t�9��9������+�-�'>�v9>-�*/RT[��߁�󄸩H�����?1œ�ˇ�����C4f�ZB���	�1�Us��"������6fѳ�yWS��D5e;h��צ����V`�jZ&ҺU���%�5藥��YZ�Mm�l��D��P��<�)�+�C[�\ ��T�-ǥ7�h���i�K�|�B�j���h�w�_����2s:']rSf��4�b�����ߏ�r�0$K-B0 =U�k�/�w�G--���'�S�篨�����K&�v��0�K��+�u���o`���L^�{�*��sV��rÞ���'ξ?���cCU}����T����e�G��aJhVN�;[	��5���~]���M���$J+U�:ϙbL4�L�Й�2��aή��	}�C����S�엜(�a8�?��sw.^S׏��8H(�"
��ڬ�n�1h�{���n0��t�mXa�q�6,-�f�R���0�чx&�]���~�H/���Sm��x��_����"�t,���_w1��t��z��]�Z�Eh"�m����Lӛ��`�a�U=���$�m-W���_�/Y�M��c��*�I����P!ij�Z�;��#>x���8�����h��B��1	.��!өd��k��W�q��سgy����R?O�X�A�=�%��䅯<�q]���˭���.e�3,�N�)���g��f�k�$�h�"��Ұ|�h��d*�E��1j2�d���vn��D���v�E�'o8��c���@U{,��ދ�o��]��vp!=�$JH��� ���PO!]�#�E���|���F����~���_&9,���a8���X],F��ȜH�����~�mv�	}|����bI�}`в�ޔ�4Wo$�Q Zi%7�O޹a:ܹ�݃DK��[oz�Zt{�nZ#�^`��h�p �<�%I����"���3T����̩<%%i�r���z��N�
I~�K�3��5�i�,��x�zY��9�Q�6��FږQ�e\�1%�d���"V�60Kܕ��=C����S�r��<��A�c����5ٮ�*�?5v"4"Fꭵ�
r�i����ޚ#нi�oL9�-~����'#���>C���a��N��a��1?�#G�an:�+:e��*��o�V���+�x�t&�sֿPp��*��-�/xp˳�a)`�p� ����j�/��<�tR����+���ߝ,����$����AÃ0����|J���moKb��eQJ��%uO��.U�a��.Bx�
%�s?��f�5�i0!!�^�.��@�y����,�زꯪ2��ڄⶸ�ɇ#
�́�J?S�f�'Ox�k
c"�C9ҢƧKS��GA����IY�Z1f��
�S6q�^�F0rc�����s;q����9���YfS	L��JZ-�
�5GQCN�"c��9�楷��>�o5��t��T?�Y�!�\5v�]m#�{\�ڨ�������U�iiή�>f�����˝�֑���[|@OҬFK��hh���E��g�y�������Y
AV�����V d�8�1�j:�F׿����F��k��ˮ�(���r��HL(]1��)�:7V�Y�����+�bhF$f�f���i��´9B(�V���DU�@�p��MR)�o{5-̛��y[��!gi�ݟ�5�It����P�	�c�\Lӂ��w��hb��!�l��=k9H�k�d��*��0a'y�TXT*A��}�OB((DBo�*�M����ʃZ`^���:_�4p� -H�%7�H�|_ucq�i��ʀ�'��A[���o�n| ��S��~�x6��$;61_c��(R�M@�K�h�E1����h�c��{���?����-���v.���}��M)�o��> ��}�Aĵ(��C3�Z��uՌv��X�>�x�VUz����E�=�/K��|�7�d'I�aˁ��D�?}�jAO--g�.��}(&��f���8�Z�$hn�p9��v�Y�,�o4c �����̅y�_�M���ZZ��%VX:�;��Ƃ�;l��-v�����Mܳquֱ0-��|��<+�.۴} �T�1"����b�Q8cr�+z<�'B.W���cd>���/+��=�ڨ�䙻�����S'me��?�=��$��*H�j������grZ#eȡ��gB��TC���
_�aqi)���ͤ�$n��'j�b!�*�?�0	64ʞ@�=.fQT�p��G�c{|��įo�yx�4m�%���b���9�x�ҝ�������ȷ]0�%~���`�T��Z(���>P�O ���^� ?u���q�>�A�g9�9�>�3݅�~N��ݕ�Z�����?���EhU�O껼(�8`̄ ��;fܥ3�!���������]���h�?	:���	���w�����F����	����k��f��@� \�������٠38�gBٜxס�Yl��<��