XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����\x�FEe?z&�[x`�z�(y�)�X���4�!��a?�����R^_���@�t>\��
����*Vzc`h�m?��^�g8䡄m��2��#�i�)�,=B�nH��;�}E�ŪC5�.:� Qy/�/�l���������5�|��
�0�����/��l�Ь���'�x�kO�nW�.¨����Mg�B�������
.(v߫͂#��Y~97F��9�5��q5���S����,�د/
!��M'E,�+�(��V�3d�v�TK��BX�dQ�l�6"�66#�Wo����r>�
�3�E!�lsy��t_[�"��z��mZ,��o�M��Ԁ��`��{��6�����u���ʺM$+�׎����T�c��׫�u/��vlÈ��C�Dw����z���
��Հ�,�	�T�ר5�N0
����aU�on� 1ժ�"��$5�@� �b��+��^����}���B!���尪$��f�U�O҂1}7���5��`ɰ�點�ᾼu�l�c�dW�կ��1sy�`�
��=,ݔx<9U�Ի��Ո�v�$�v%�!8�n���x�:d��2���7t��0v���q�Jk��T���n$�墊�u��L��-ؽ�)kxg F�I�W�V�e]o2��Z)Yq�=��|_<f�P���ptƷ�q4��&���ЦI^Uf<w%��JµA���:��}���q0�I��Tu��.��y��գ~�V�d����P�It'�q�[TXlxVHYEB    48e3     e007���*2y����q���[����ЭFP��%f��j@��GE<r��f[~��$6�G�U�M������#. ѡ�pI��]�����0="�X�b�>Ǖ`WBDc��f��Y����9Ĩ%Ȟ����{�{���F�n���Hzn���w�qu�_�Hq�˼G��n�hz��s���EcS�R`h�N+9�W���R���o��YkA�i���O�t���hA֑����:�N�W�S8��ل��>S���F��:7o8���_�\ߴ��!6w�ۢosĐI��ǝ�1eB�q/�q�:J~�2ޑ��`��f#��.��9�su��b3Lr8_��l�΀�vWj�a~w���_@��w��0���G�^UyA��B���H���e�U��6��*�jZÝn4nnv�.�T�߁e����� �o�ڂ�,?ʕ8�;�����{`{�ed���/,뽹6�c���N1]�In���� �(KC�i�ZZ�G{Ki,�d��;jѿ����\７����f��;���o��v�Zڐ�}\�nr��C��|�8D���Ių��wĂz m� y���M�,u���os����`f��ma,��f��_�ķ�Z؀�<�Ư@0���x�ЭQ� [����?!�s�zگ>��]Ϭ~�V�N�M\T�㔆C�/m�� ����`��$
r{�<]�W�P{�x��)/k��|o�،��Ƶ��.�6�;�䬽�H���4)CMdȬk�l�/;��y,a�J�<� ���[Nitxѭ !�U�!,��L!�7%�ޙ[�wɨ��ف�W,�4�x��<&����搨R����f_�*�����\��w%��:Q`�F��E`D��������=�Pq� �r7g�O*q�PN��e��\�Po`i�g������YC����W~����Z�h؀�ZHY�G0So���J&�V��;ԆrM�������nr�����xB7�S�����G�r����	`Ơ*S5�+���2ws���4L��F�s���T[X}��	���s��3�pڷ����)+�\�N�[��}¾i荣F���[
�k��L$tc'r`�'���-�Vܐxj���CS^`_F}��&+qȋ ���e݇�}A���,'N�Ac��2 ���8�`{�2oޥ¨����^�Ү,QĹE�#��R�S^�:��nN�-tv�]�;���_k��$2ut�E�em�R|r_���d�d��g$�1+�w4�F�2}��zl;t]n�g�H4.��Qt��H�I��4�Ѓ;\
�d�?�C�1�K_1q.$'���V+Z7/K%�NA[���/��e�l?���wi�������#�V�2\ .4	�Rz�)��[`/�(��#7��g����3�j�N�H�t"�p%��r����q�C��3���m��z2���]�"��ɮ�K�o�(9Ћ��7ab���� �1e�#�����%��*��nW��������S}(�`?��3�؁er(ϕT����1RL���ھul�j��a{�XY������]V(#������B�R�G��0BP������a�V� �l#جs��Q�������*|���S�5T�,����2p�,�t�fX9!�A�2�Ĭ����c��:�����:��6<�q��@�٥�wOy}!��s���(�n�d�2 ?ʐ�Q;}���?���P�*x�$P��U�z]v��$|�����"�B��������s4f�f"�3|?���_�L*�A߾hi_m>D9sj��ka�`�k�����K��
�����Sl������o����
]uPTj�Pq���-BEGW0���q�	0=D��.���wm�(8V~`��Ԃ����x+��MR��XO��>�ڏ|�r�3��4��,�I��Q�	�����2 eO۸�j�����L3���#��x�D��}0�Ezp�C����B�ԁBe�&�l��.I���dc	ڬE��<���e�Z�"E�{�L��Z�G,K�GȈ�{ۖs�f�l�ո�L�<����K�ֿ���S���:'�z뼦M mc�O����ub���.y� &��`��1��y�if���ܱ
�ݬ���bJ�!�t���bn�w�˼�S����	���3���bPLj岯��&�ɭѮ��u���`��cEqu3sJ�ZKF[����Ĺ����l��:5U�QC`�Y"��8����#&�9�Nqu	��\�c5�ӎ�q�	+ ��7Y�UGC����7������5��MP?tC/{nF15�r�$�8D�/�J[l�0-odV��z�s;����#̍��A�ҕ���*���!܇�O���
d�6m�23q�clQ>p�I���|��lB��h��pT��0E �+���B�5�v�l��bPH���J���[�la�5�HTE����T��-����	��7��Mtj�<'��@$���,=�|��{���#�.-�k�N݈h���&y��F䪰Քd�����;�3^dȌ��#>Z�#��g\@��	�*�"e�7�40���sMX@�"�<m�*�>���r�������P/!�B��z��g� |�G�i]?`Qe�wt���jo$���*�������m"CL���������p�iO �`�����sh��)&ln�`�LU6��E�3~>;���F��*�}+�Fl.�x��u�R���KKbw���M���T���(�	�8[�z3�>I����aM��ȹ�mEl���J�Pg4c6�5?�y�Y����Qym��U�͖��ni�-��/ȝ�z��4��uŐ��Fv������!,�L��w�;�b�pgJ-�l$@�[�Yy�m\5�$�#�� �U���|�������c�0"���e�*�,?����� f�*�X�m����U�پ'���m�YfUQ��V|s��*>��VY�w��8��{���r�Ni�d��e�1����Ɔ��퉏$��*��3�!m�h�/����C`�F�lςF�8���x����?
}i`)X'�iutƷ���9��m8���*[���}d3��:���jj�!���Z���v[�ߢm�X ��;G�� �a�QÏ��L89�(�`8��"5/�b�q�m�	��ſH�$��+T��Q%���"���x��"}�Θ�"�b��q�8��[��`�FB"�����Y?9�Ⱦ�b(����U�0��$�6U~q���s*e�v�ƹ.)\{T�d��X�����ǜ�`�,?�r����iͅ��?��R|�i�eͯd��:$��^�=>��P{C�h��	�J�ѹe�.+ۨ���������z��Ķi��E��ҫ$�+�"ͽÜ���Q��-���G����t(��/l��y��4����"�[��&ޙ�[�yEs��<���.}I��	A�dv��t����U5�]@�e2"�/���Uk���ns��T��;��SO��� _#��7�o�^5^��Xd)��X�'��8��4H"��j��]��#��� W蛈Ig