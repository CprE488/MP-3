XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����G1+�.�qr�{�~$SΥF�����C��$���ɨL�mC�Š�B���	�J����u�-�:��¼��c8�/(�E�� ���w-7�Cfn�yL��sJd�ϵ���6���0qߧ�E�4("�R7I���Pk��rfw���Ps${�Lpy��i�M
��IMp�`*��f��27���_�&4��w���m	m�#�'���L�~%k�EH1֯ꮭ�-'Y�2�S�$�����nb�w���Fx0ı2s�~I_�s�����V���U�F�������Ir�<ħy�=�^�_{�O$Q7�8;
���R7[�1��~����X��Vu0 V��^��Ւ���s��S+bt}3����j����X-���\G�2c ���N�7���=xp���&�+��#2���R�m�1:]A7�U��΅l-�+�7���ƌ�ON�W�nj�"�O��mk��°ך�LL�9��/��8;�<�������kW)�G�m��_�o_E2�q4ꦿ�n�n�%��3����T�;$��\ͮV.m[��B���/�?@�s�F�9�.�Z@��	���E_�$tӡ�I�f����f�K4����C�̑��wZo�r��� ,�\��ߊ��m�Vx$\���ȗ3� �����j�{#;��&6�A0�t���'�'�H��
�s[j��ݕ�a\��C	���8q�8QN��W*��ɾ �o��,?k!GKe�'��W�8B�Yǩ!q}����1�����D��-��4f�NXlxVHYEB    9fc7    1fd0i�(j%L�g���Y�߿��&�t������p�p�?X66Sld�Ip�h��+�݊�e�ƩK!^�a��8J�@L[�>��4��=�^������`D���]������rj���ʋ̐�ځ&�)\d�o
����4ގ��C�7�����8�b�,Q�+��K��}�?��/l����m��U��I;��n���*M�"��u��v����c����p�|�w����R��.� "�)9�s�_(�=��'��41��5e���CF'�|�״ӣ ��wN=w�[���`5=qL	�,�k��i$m;ײ��l��z!IR�u��;3��&.���g8�K~R ��,�I���Ol�\.toD��o���9�栤���/BkM#���/j��q�;&�ew�9r �pq���*p��[9�l+��B(��8Tl��m�S3;�Uߗ2E=�k0" �i�.�����-���n0�o���(�T����ȟt�����?թ`l>ߥZDꠧ��<H�YR���IK6��/Y/`D���Q#�;�;v�i1�ÊAG'�M�4YiQ�)\$�K����LO��3����O@{��@X�a ��~#&�zY[�?�6��nh�*�P�J�	���`W�p�Jٔ[��ݣ�Y�N�0����]��/Z۟%cQ�рd#x����#� :.v1�C`A�r�o���^��O�Ix��"u�O���Ȅ��{ �ã�/ٍ�lV3p���U�&>1�%�/�u6��.A�S�H�Q4�`P�N�z>���LÌEYCBV���㖐zl��j`�-W�M��g7=B�S��Ӧq<l_�酯�8�OxW�&Wrnw- �^�y_;0��8���%?�P�hR��Byܤ\�E��p���a���B�zkbtx8���aIO�4��|��M�}S*�������S�U3jÞ�&��7H�*� ��b-�����<��˧�g�yb��qp4�J��4{s�c���C��7!
"ԙ	�D�G0]hwJ]�|(��Y�� �	�׿��j���Yɮ���:��@Vn�u3(���>�)*F����B�%�p��&��"��j��ש�����`
1S���O�?#��*�ޠ��A	֡�Ig��˿�)�g#�g��k � 8�6������fVwFHA;���=ML�g~���
h{Iw��D�j�G�����4����)l-j3r�)�H�h9
R��&6K�S���G�k�r@���i���E��rտBX��Pw�Y��EO��P|�u�D�T�
+a�/�)t�NA����n�6����t;NbK���`�p�PX�bA�Η>XI����zŰ�msX4�~f��#�l��Y�(Y� ν;P׫��������W?@fNHk�M���-w�2�Z�ӓ�BY������U�J[��O����4w,W��E��C=+��~�|l3uu.WOE@���0f�ાs=��I����C�oj����{����4��P�(7�bc|;~����ޗ���)���!�9��?�o
�L��%v��J�����]�L @@��Cl��XR��H�f�~^͋��u<aM{��Z"��X��湀�?0W��W	>��JQb~���WU�#� *���:��<�:�'`�*����oJ֩�7���^o'��`����=Q���O��R�#��?�:4�$��n�$+�bd���k�,Ȝ�bf�/�{��n���$.�\�[�=2� $~��%����ԵϢu�Ɗ	
��^�Ow����/0�Bw@�Ut��C��|`8�J�@ceSe3�;�O�g=��q��r�O�(pj�օ��AYHv�2ލKW�Z^Fq�A�t����h�L�؆���Xe�C��ǯѝ������a�%��-|����I������U��B��D������v��v�ں#aT�v$�f�Hh�b���My�f�;�͛��>"�9��J)j=ɣ��h�����K�a�u;K���FL��U('׵���=Aܕ��KOe7���F7�5�M�R~\e΂�Y��Z��U��띘�Ւ�{���(lnO�(��Is��k'*E��7���D��by M�$������~�;�a�Wo~o��ݻh��:nU�� 2����W �/$�p���d'mﰩ&�?���3L�Ÿ���e�!)��M:�J)�v�����'���J���eP6&�S1*���?��pd�ă��)�;�CK�ӟ����E�~�qj3e+��Ճgƙ c���'P�i���[l�	'�g�/ͺQ3�D3��W�L����(��Ц�r��Ү�p�Mm=���)X#� ȑ����Ti������A�������i?=�^&��F���ic���������?l7�w�����3F�(�y�~:6�Z��RO�֡N
[������Q!���`��?��ﮇ/��.�/x,Ny�b��?[��] �^�RϩR��^�gP>����a�l7�x�[�Z���:e� ��9*����1W
Ӗp�=����B�@׽�n�`�v)�%�'�����>?�+�D����]��`=Ź���E_)�y8T��C��J�R�v�{����'n����-Y��{���Y���[�k!'=�ҍ~%��D����HY���Z=R�2��y��l9|�~�\�9U�E\ࠐF�tt>K��hC���rl�2J}�cU�1��c��U7��&�S�~�H��նq��R<��6�δN/���)Ջ1����=�c������d���i���H����M�'�.(5I�ľ�3ݦ���HϓC] �j��`0�bW!&���%��%�IS}�b\����� oP�2F,W�,�8�f/�Q�����A��!�ڪ�Mj~��\��	a�JbTH~rw��H�FMy#5�Z�x�S��,��� �������;��)��(����CP�b�W��x�v����X�ng���:�S{�|4�p`н���S5��:�g�j'���JP-�|o�_y�u댽�������Z5�.��9� x��wk��$+xU"߳�Mq�kJRw0�e�s��d ҷ�g*vg�4��قO�m�6���y�#�Q�/�Z��U�`��=bb0�H�%��7�;!��\����î�ri�[hʁ�؟_�vL�e��\rJ!!�y���&�i��m;|� D�=/�^�� ����#�{����,��
+R�gX���E�M��5(+~���'�m/ok�>�d���$)���������KJK����R��[�̏��/n�@���/��䠹:o�C�0�T_� ���/�aB�j�=��c㸩4�˩���Ï�qTS�����A5�Y��LF$�B�r
�/��=x�cq9,<_�Y)� $� K��z����E����ai�������>�j�-n�f(��02�b��-NK,��o�y�֨�+S�b��v�6B�A��hHj/��@��c��v�Y^.`��}�c[7�?La+��]%sғ<�-�Rk�H�+ic}�R	�6#��gr���
��e��~~{��_��;��f�ί���wc�U�!�� /Ƚ�X>.��2��)�c��D�Nq���������)Y�hh�+�������snp
���:����R�����6;�)�p	 �`k��<I	�l��I�'��QA�w�;��9ד�P�3s_��$���<=5ږ�x��#,�H0�/z�ym�j[�h��J�����\w��]��ֶS��E�>,Ȅ�+��pXXw�n:��שo� ���J���U�;̉�$�]�U)f��FO�;����ln�԰��L���c�[m�xY���3�1�.���ֲ�!�-Ckպ�z��
���-��q�s6J9�E�ٝ�_���%s�k�S�ݸ�t/��W������Sa�4D�� �^����T�0���e��*j���رl��#ۄ�I�����wV6@��v�;p=Y��&gm���q�%��Rߘ�^ߖ��^T�xu��sR��e$���,�p��%�"RhTk�����W{�t"}qh��;E����g��h,�Gc��� 2��6�zy��	��[�\��ۏ�^	Y�G��'�[�ؿ��`��J������6ߖ\\��zK�U=P�dҶ�M���"nz��QH�-b���'l�4�.F�jv�u�J����n<J�ۿ���ϗ�h�kds[�A����>�u�+��h�zj��pV�U��ϭӯ�2���e	�m�^2B��[x	�E����!��׋*�� 3!��8����ν,y�(WG���\�=��8��x��p��z���s'��T[�ܭ�L��O�27�����3��a��!o�I�=ᦗL7h9�m[�ܡS	�ˢ<13r�ۍ~�����C���+;�����l���J�� �}�Yt*=(H�X9�Seկ.�VBP��~�
�v?W#����a枈MPU~g�E�T8r�0�cg�	�xݶ!S����g��VV���AI�Nu_)��gK�fa>�N�a�H#��ҩ��97���^e������c�C�b�]�~���J��;��^�J%jW�C���Z��W����X�4<�#�Ծo?wK�Rc6_i��V�R��lk1�Иف�D��.5����ڙ�y�#~�W�_. �y)=���E:�=�O���Ӎ�e��2!��hC��?,�2ZfȄ�n>�.i0�����G�1�S�=\�T�R��\iO�XM�4o5�ƫuo�x��5X�
�O+u���Io��1�u㸚��.�Va9��j.�T�m�!!��o�I��Jf7�+���:9�s!^�n*ʂ�U�,�%�eE�<����wd+Xv����"�"{�J)�ڿ(��$ݟflQ�ں�.���A!>�4�1����n��%����=o4]ɿ�3>zf�����h��\�o(ӱ#������y�_,).�xN�໿Ε�xF�[�������՘�(���h2�ݨ 1g��an��^�*;I�B����� ��~�HNW�6��!���+j��d 3��ج�M��o9|*�0�2�߻�M�J���R�0����ըP=� �0�d�z�[�`:u��T?rC�˝����m!�\a���6B��к%�_j�D)�h���\�;�}�څ+�' RU;��w��-��(�YS��vh�6�����T��z�����a��se�ŧ�ӄ���x����J����`~(i��#����B�bLW�>f8!��n1���{��'��ȱ�K�����^���8]�!>F�Br���
���ռ.��K��U��U��o��ډ(mb���s]}�.�,F�[��0 ��$Y��G�e���o%�a�Zc	O
�2�a�^�\�Ru��`0���{j�K~?�i�sS:�Ԁ�`���pQ� ���gB4rі�5
�򌖖0�Z�q`
��+�,��NN/^05��W��sH5�3�Oa�Ŝ']#!g~\�"��s
,H�f�2?��{��	�U_�$p���.��g(}@����!�D���b"k���돶�A?�O����m� 5"-N].��)�e�� ���6�. ���B���p$�5��/�C�Q���7�lNUo���O.�}�z��sF�l��9(���'@1��p����'[��G^��M]�}1�S82��Rw��<�Q�p���B|�$xE'/-���l�N�ώpI�Q�����ot��+�s�(�k6�9���!l�_ޱ�	E��LBp}p��
ȵ�������@��@?�{�4�yW�EK�|U����I0?�6F�_�b��C��<�������e)+�BE�Y�:�$*�E���c^%��_k�0Nb� �hB �f_6,_Q�7��k�qƒ=��'�t�8k�6@-����G����A�9ElNqN&R��:�u^ڟv�oy��d4�D��'�ӓ`F	�r�P_��Q#B�V������I+�>����e���RH�[�wyJ�q�w�:����VS��e�H(@�Sg��b �A�k�n�S���pj�n@�R�_�*�"mj�H��5}aSc����t>�r%=�������~�M��&zsb$q�Ӧx�1u���p_`��B&���[����+�c2�P�J�4�ҨB�r��N�ب|D���Kձ��!��O��7+>'�?����:�ޚ8= f�:���@�O������J� �gc"~���NÅ��uN�;� ����;�RX�.Zf��[aAz%���El��nS�1�@��/�t��T�1����L��S�<jĤ;��f=�/�t��L�)�6&.����0QS�6e���1��>��dƊي66Y �*�K���yLM3�u�O��-����g
O52i��#3܁F�Sl��n
Qi����R	�2�(�f����|_=�����ֶ3G�Q$V�܅)-1�	;��Y� EȢ����m��4��f���Y<�u�Df��� ��hxoY�����[�9'0�Mg�W��.����,)����S�i{>5�]�d>0�IA0-8�="k)˂ L�����]��2٨l�P2�/�S��2��BPg�,s�A�Cq�y�j��0k5�~S��Hb_@k1�x_	����Ǩ�{ker�ڹe�M۸����.Sl���b�aq�V׷B'���}z5��h�ǂ�K����L����O�ph���X�}���K��F�Kno�l���^Jp��o�!�3�
3����y̍��/���[�,"D��| CI����}��
��Љb�-��� >���=iԼy3�h������j�[o�Y�<Ư9�_�'��#�u���V#�*�X~U���}����r�X��/���SȺ��1�y����w@���Xw�8x�YӺ�қg�y�6ٰ�Vpg�	�Rݠ�@%qGT�s	iH�ѻӷ��9B�;�/.�׊��?���=-ʤZ	:�+�:Xhű?p!/�Ѵ����ͽ��!g�I�B?�f�M�Oo��6?��L��:l8#�@C}�A���Xu�Me���L[��Dn��NRe�Ʈ�n`��||`�1fu��V�A��`����aj�|3"�	Q�����0~[�Y۸PK������/)��˼����i/�r���ޒ�Y,��䍐jδ��s�ɳ�Q�����=�U�CU�6����f��1�T�&J\����ZRK����!lC$p��䷱[Z��O��7��\j5���xT~|��� 2�g��a�goE�l��F]�?�IP�"���؇���1��m�ӌU_�6�J�/;J�@M
�������>!��چ^&�o�l��| �;!��Q�L��Y��/))&5��N�J�g��f@��х꬟�s��v���}h��)&܊���N���H���D]匛6u�	j-X�1?�;��Y,J �
�-C�.�6�/dϻ��A��� ?8���Z��]~el{��-��8T�{h�t�t��m��Ȼ�(=��70��6\ĩ�S2��(  3Ig�@ ��'a7����G(�"��@ jH�OrJg��b�yPa�`U$�#��^���!@g�l��6�5~�a���+��R<e���h��q��|np~c��͵����
j����č��[��]��g~N�>~�A�7�a�����0�_���N�����|�����k/��5���jG������#����~�ך�� �%4��8㰸�H(��Y��C�E�Ov�]z�����Rytdw���'QH�����0i�>V��ɨY������C*%M���M�V�܊��*f����/��#�Ў�҅W1�L�����Pr�w��Ȣv~�TL̈́=d�+1�J�F*��51.�n�z��
��eQ��ʂR��^��	F��5��1@5V���,�>d���t="w���֦�D�d9w�Y,R\�ӕR��?xF�`l<�!�S����j}}S�޷ܻ�!��W]`R���J��_&Rq.�O������fʋ�;щ�n���y�C"vY���ʹ����ʥmݓ�_ZdË���q��