XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���R݇���
(�#���T@�2ʸheY[�o\�A�����*�Ll����q`�,����w�əɍ��af��A��W���B(ٹ5��ы��Q.j+&0�ݫ
�j�SRC�3A�0N��QU������'�Gr�.q��Z;��s�$���z��`پ�ݢ=�q�ڧ2��e~d���X6�l�Ն��Ƴ����^��17?y>��?���EnuF(���(��4�d�3�W%_���Vx8�<ި��^|��q@��4>ӝ��_�����BX��Q�ڧ�<Ϻv����ܞ��	��Bq��l�˝@�UY����E�T�0S��V� p��y��D�ə�M��>��u�z���\S�(&׹*���E~�]�/�b���Щd��RO�C�_y5�C]t�e����S!��@�^~=x��:ۖ�t�@.e�5�
a��v=�=I5;��e�A�Gy�<��M���J� �;m<�@���ig;>a����k%4b4L�z[�'�/�1�M��IN�+�H����fC"M���]�s�g��ƚc���H�F$�`�$�����X����a� �n}�r"�"�H���N8��}���2gWqi�i$�X�H= ;�x���S� ğ�Ё���L��:Y�WQ���Q	��"�Z�Hc��z� ����2������F��{ϋ!Ƴ�Y<�FMpa�@����_�T�/��Q�EKf��Dx�x,Ml'"U�³�8OW��>$�����󄦠��XlxVHYEB    dd8f    2160w0�W��&�4�^el�	͵4i�]�� �8D�X|<}��7��&J��ɽ��C��-	�NCS���u��Z���2��#��"p"�k��r�gGID���3�`�	�H�䄅�b�|��o���RZ�f��KA�?K���z�,�}����f�7�'<�G��#X�����R��2�t�r1�X��K(?���@/� `F���sa|6�SI�bM�4	�J�8@��I[�:Q�%�]�mƼڦ�gF��W.bkA\__32*B�q�#Y�ܖKw�Rk-����UW�f=������#V�/���R�L������}(e�@��h,��U���@T��/�p�D�yUYR��}�3��Q0�S�&�f�'R|��Ư��y�(��}=ͭ�˶߆��m�0��i�ac���iSs*Y6^t��86=�bw.y'X}����J�5ˈrx�]���yQ�������6��Z��T����p�.�zq������y��5XV�z��z�	9d&ҮZ�klاLYR�._^u��M��f�!�Q+W��s��)+����h�6pC{s�ZQ��h9������%��*h=��5�?^$F�Cp�u���@l8#H�C9��:�]-H��\B禪4�#�E虄t��Zz&��j���@��ؘm�(J��cb6�}$"�<7�x
���n:��&ӜRn{8���ź-ܤwRw�!�B�l����2Ъy���#�-��ߖ}×���S�RE����Ҙ֪��1�¸�t�Y��HT��y@ߌ�<<7�+{��U���57ѯ�h|r{�z�vkB���H��~��i��=�Z���-u}S�����]؜Q���c j�r�n��:D�}��,��1W����Ҝ�_>���n�Q����Py��[�h�鱜"ko�bO�5T'�:�u���3�`sB��ץ*��& @�D0�#�d��%5�=Y�l�e��-�MՉ�O��D潓���)���p�(�����%��/��A؟۰��V=�Օ��Tl�����֎à�6��N�ے��E�����SfN�J���� �<��������r)B�@O��$���[6�����؁eb4�c��ijEج�.v�V���x<$O�M�������c\*jL3 �a���,Ōq��Wwn�{�|}��J++ G��Y��^k\������z7��w �O�&�d�Î$q�*�W�Ct_Y�Vw�o��x��k��e��4_��Z =��b���P�잚Wke�$P�$3F���zo�˛K��Oג�/���a�9���f�[��L���uH��Qz�����a��Z��x���m`ů�4��yU��%�
5��m�-x钄�:(j���(j�p^u�����AC��w?9���"�����ӡ0=p/�k�;3p��hҹ�.����W�Whm�l��l3�_*]��ޕ���y*����`�9ړi^���U2��(f�5�# ��,m�\�|��}UK�}��c���y�`��y;m�OM��M������P�r&�צ`F�T�n"XLD���%�Y�]�m$&�\���B��9ߍm�3��G�w�ۜ�WH\\�1�h �/
(E�������7�#��m���0�ay �P3�Nv��)`�67���=�_��3'E?�xs���y�L�[����g[M6�Ҕ"7�㹇+���9�y�Z�L�v�7�,ϮS�����EH��}L��>�o �L�/!��:2��w�8�N�����d*�4BXhG�������n`ogŚ�����[x�8�)���Wd4�2p��A$�۔1�c�T.�Β�� 0�e��볢&6`��f)_��c���J>2�A�BeA�y\�Q"3J��~�C���S�����bDfx���+A���-K�0���[۰���N�� ��811�5�!~�$�i���j��X	���1.ڡg����&��,&�?Ujy��(�^6�����sw(��sR��3 ��̳������(+Fc���ʧ\7�k��N��|���}��Gi9ɰ�{uOوig�7�@34� )
,���%�S�/��]G�C�X��vK��|�sq5t���I���Z�!����yLmݠ������rZ�:��H�/�J�����fnLh���8q# E啪3i�5��2SR��W��^�:�y��Z6M;�#~Z�Px��`��Л��[�ze��S�GF��2M�m)���=-z�~�eT%��R�e�3 ���%�B:/ ��8�Ť�����)�I|&\V�|OTh�)��dWU/�p���|{�:;
x�2�8���I�Y��Y��.-��
n��+��"�S���rr�٨��r��xE��h�� ��+��(�5�E��D�Z�!��o�Y����rɅQ�z�f��i������9*���ȝ�B�$m�bN�}��0^�#������} ��b�'a;�-�`6}��I��}���L�R��N�o/�����X_'�ۏi@��N�蕍8O�1{�`�}���%�y�C#*p�]���`$�3v����x�U�;z"-`�ǩq�U���-@ �y�9n����F��ȴ
�Qu@D�H�-�] �^|���c��1�|�-�g%��A�1����a��U.�T��7��M��d�o�)�9+%����Ό�:7 ��S��rB���o�*�Ap��KnL\|(��x<#`Qo�L��fr	,#3p5- �6�KQ��Bu��+�z.�������G	�/�"���z���_���k���ٯ����!2��(7��X�(e��e�
�j�ok�������<T�C@����҇Sh��fE\��U��R���k�У���M$H��lx�@�0pq^A��*t�����Z���z�f��*6~xD>�ę��iV���~^�\��l����`{&!������,�s����e�a��*�?�߹���?�i5���ED��k�_�0Mΰ�D��oV~VPM��B�*P�����g���h�]���rm��a�h�l/��ۖ$�-Fi_o��y�������#�����d��\����K�=ľ1�h0��p�úN����7�΢Y���bD����O�j9��I٢
Snl���N��y�㲖����A��g�xd!� B�G���IJ
(~�Su#�5���� Dˑ}ws��@'f��t����@���,8�ɪ�i)rۧ��]��;_tU���U��A�h �)�����1����̂�'�k��;�T��h긔$����<
"@�8�E��5���x�R����Ո�`h���ۻ�GIT�&�A?!��d��U�Szt($a�Qg��胬� ��ѡw�	#�łG�3�` $�IE#�3�}��#*4|Ү�n�k#0[`oǯiD�vБ�@�/G������d�
Z��=7LW��)Q�`�+
,��p^{]�p�<���оZ?1�Xa�[ߑT�����/�:�)働{y7��7��r苻�O�s$;�M;?�Q9>��Ѥ���%?��K?N6�Оb,�1Đ9~ᚭIc�X2� ��H�%sF�!�1@5�ܜ�X1�LS?OIW��)��=ٴߓ�����@��-���c@��$=,��eݘ�Sy�;iJ1�OoqV�Ƥ�qYw�U�ڋ�O���|���f�|�S*����<!n�|��_����	"K;+���@��ڦ)����"�;2�+�I�x���@�N��&;\zc��L��Cq(n�l)c:.��<<�c��l�X��v��R�A�]�H�ϙ����C�7�{o� 2Q�z��ۯB4�@��k1c>u��������:]s)P���;ه��:���l�fI�|e�"��P��ͫs����?�1i�O��U7i�P�?�m�
��?��VNJV�u��<�p{�e�����д[mL�b��<��4|�����@q�~A�d����q$4]2�jM.��H2;��S��f�[A&­��� f�&N���5�#T�m�d�{�ۋ ��0s���'}��>�D�3�)��|��s��fN���qfcjo��rJm����ҥ��iBc@��+E�����^��.�� bA��P��ߖ�8�%�a�J"D�� M���ܻJ��#� �) �S�d�C4��'�k���,5���z�~����.���x�a�O��`��CI���1'R��˗�GB��z�aІ_$�D~:���0/�qzr�rU�I0�_x��_���4hu�����3o����r�	TT�f��]��٬H����G�`:r�K)�WY0�*�p��b|��Wu���și$�E��IU�ξ�����@�����Wj�SG��{�o\u��W�r�;��lh�[��:��n̩���C�Y����:<�6�����	�" 娵'�#���\���%��%�f� �Ԙ��� ة���ul]��v[�)^�,��^,&1�)?y4�ᇮ�*Tz���c�����\��E��@���	��t�۶-��9Z:���duvqG�� ZB�p6�k��
��{ߒu<N�й9��~:�MB}[�_��������뷍��������J��O;��0K������$�
y����^���-�:��b�E{�%�	xm��^��$�F��HJ��d�h��Lz_P��@P��6²��u^�����r��9M-��J�I�<(��^p������W��'t`���aa*�8�7���ͱ��Wy�L���QP�rx��gΐ�o�ߢX�{vm���A����Ě�VF���6�9%j��qٖ���4>���<�5�A;����`��9q���n���D���eM�{�跩��	pe�{�R�B�F�03�.�/��/8ͳ�fxy��������m���o;����Xt��y�,�v���ʏ�䄉���`M(��#��ϢS����N�g�x�7�2"���f[m�P�»6 �`�,����]�J��d�u���:�f��?W�s&q��	�>�{�5�m�x"�'Տ�z��L��8�����?g⟤�wxG�:I�}��ۦu[�K�{�h�O|U��X�ʤk{J���8�N=�}��'Ӂ⥀W��:���br��cZ@�[�Ϥ
,�_3��r,��5d/���uo�2��R��q�|\��UN��A�������bW�oxIq/��6�ȟ��ׯ����Y�Z{�B�YF��%���($&��0��Q����iE�Vk������rl]����t\峲*۪� Q���V�����A�m��Ų_�;���L����umF���:�n�Ҡ٥7�	��&�����
����A�3�QjS�6��gд�����u=�j�aU�n	D<"��$Y�X�PDI�ݱggC$�>.�y�W=�H�s���-Im��F����;�R�hB�-�f7T�w�_-��(1�*Tb�~]�|TΏ���i.YV�pAI[n�:0���ΰ×,I�]��~_qT����}Dn%o��\����7iwtK�ˮƅ3�����������>)f*�(k���X�@F6/T%8��X[A�-��X(�@�-�:�U7d�:��TP��j�q�hU����>~����P2Z<1�?KA�v�����[*.o�@,Xs�W�F P�m<o�F�*�ʑ�=��e���<��vč��P�GE�. �	Z�YA�+8Z��:��g����SD��ڨ��:w�/7�QW>B0	��>���F,z7Y�tc���w�7���*%��=g~AS�ڥ$}�eHͬ���9���M����P������+ �*���<��_�NߨYGFT� �^s�V��xKS�[H�F��V�S�U�ct�2�X[b
��(
����l#<(1�z�v>>��5�;
p<U�E��q�{*+ip�L�;���������ځ:$8��Z���!�C���y0׏q�U���a�x�AJQ��V�Si����D���vkhU:��t�DdK��'x��*��Ý�"�L���c�V�$��ļ&���Yɍd��nÎPk۷�@D٧��DIX�P�"eԴ"��U�r�H�@�޹��Pyԅ�n�����\W����d+��Dɸ��������	Ƹ�F�+�w�"�5�?`GK6�^L�ܷW��������1?	ʞ~��bB����43����姙$|4%��`dKm�:	��g ����Uq�$��T���KQj�sU�����,�6�q��.�������H����7a��{r緮�/?���>kB��'���\�8���[�B��_�^��πf�|d��$�o�}Q?�}N,�Sq��/w\z����q�5�������Gq�Y(���
�{�l�UWk�5h��r��:�RP��R�W�Hz�w?s��ߡ���pӀ5�*�7+�?ʍ��������ǪD��L�nk����-�&����Ժ�Gv�x��*�!���/��^�4~�-^zp]�����Dٔ���&������OX�Ҙ��OX:FݖʒI���c��X�'>�A!��[9�&z�#t��a��t��{�1�Ia���a����(�m+�%Ђv[[���8i�{��sA�����k�(��Җ1���bG"��0���Q�F����������m����!��Er18����`j⵾1Sbsd՟���	�l�wl>s��:;׮�1�l���6�^�4��I"�b�h18�쏙�����A����r��+0��Yń �/�wH|�+���:	ͧҹ2�\�_��|V1�Y4�i�yQS�����_�R%�J�Nˆ1F̀ԑ+.ûk�C�oQ�%�F� @Cxگ���k��	h85�s��;&o@�z��y2l�;޺�g�[L�j�c*�,��UT	Ӎ�ygt�T.״�Ô[���hjr.t��tЋي|0�1������]l� %I�w�l<"{zQ��uڵ��,R����a�G2��P]�;�8,	܁�_�V��̡E��$����+���{��3����{�,��*
0ڜ5!xE�h�]��bEM�R�f��~�'������F�@F��^2�L�`T`@e��8Y����{I���"ҚA�9/���$���1qDȾ���J�W��=u���� {@����qV/tȻ��f��5d;�����,��ȴ���N$y������bX��5��o�v�y�n�F���F����"-�	W�BA)LLN����`h�8ݏ��GPբ�ɓh���מ�����r"��!�ڐH���֕٘)��)Ŏ���4C�!\�Kol?ʹ���=ڄ�Wl�����
Q����*[�V�ڴW�gog/JlU�f~�v�K�d}�G�	�z�ȯ�֧.Ι�<u;��.��u|��ґ?�h��ſf��@�k�B�W��v�X��
 �F �?��������ŀ���mCU;��w��QE�����`���0��w��v��̑�h��U	�m�N6r�ʢˌ(a����ZTL�?�'gۃLX"�g�:Y�-��JeCӢӔW������p��:��]���)r��VEn[jy%�Ou�$AWz���u+?�=��D��> �^��Ζ`����<��BGu ^7�/�t�����<Ng�HB"�C/I�������VbA+h�l�su�ZC~wr�rQwh��XpNTt��`�+��1�Q�6��kTr9����+B:�tq��FHm�mv�c��:X��!f���f��ኛGy�SU���̚ʒ�~���P��vp���e�G�9��M3;�(���T�$�JhN
��w���R�RQYqSs��A����J�d�xM��F����X�q�Vc4 ��|�Q�2R��W���a�Z���1�-L�%-�I�	@I�eXK�
�(j[��;(ُꤲ=����;���w��M+�ʪ���g�g�x��b�Ј�ذ�O��e��>��ݖ��Z���Kˋ�W�E�(v���LU���?c}������|���W����P�R
�`�ٿ����hm�{G�}��_��,��G��#�_�
@;4 |�O쇌L0rߩ?�Z�I�/�m���.����?����:hދF�	q��+[�6j�Ȯ��w�9:��,8��ޗ��-P׆l��N��2���z)I�p�ò��8���8�;%�膊@�|)�;�s�;i���$�kÎ���T�~��_��!ي-��V5�����t�t�d�k�R����-�~�����h����
�X��jq��s�X��`�+�\?ZK��w�1�L����>�w�vs�'�~0o���U	�h�虏ٯ��7��+��h��������������uE���$6{��X�6�+��~��(w�N)��?qud/g�)���!Nɶ��w�:o��>�����>�����}6!�HW��