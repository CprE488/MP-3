XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������r�Z�/ύ5�YGBKІ/k���١��Y��Y�6��ڇf�A���4��]���(�=��\���I�W��N��}��	\��	g����Y"�H�6��*e���D��AFT��ߥ�Pdi��y�$�M0���x�Ƣ���t�3��'B��n�Ì�l����%FL�2]�,hq�ǀ��7ep�n�E����u�,zȠJ)^�ǖ�� "R�U��I���\��C\�U"��r��^O�zc'Σ��`q��9̋N�S�go"���z�:Z�����ɑ
�������gp�E�(C:�#e�#��Hm٭tZ��|��u��ϊBݷ�]�ěCܯV�֐� Gfc�����g�r1��q��2�B)��_�7V1��^y!�?NLr��`/g�G�B��(�q�I��:@g���3������5��7�Ͱ����|�+Xȫ�c�-oQ��?� �����+�u% �O���E����r��_[Fƞ�q�`�8K�\���{��02�&��R3�QO��-�^��u�kӂn� EV?�QBIG-X���N��+���F�N����B��>҇!�� �J����!���w�߀K�x;���p��	_5����'@;c�D�Վ
dbp���\���p2=ab��*���A�A[\�;���Bs��ken�{���X�+!J�ėG���"���o�O�zV��y5|��J���YZ�RXj�'mf=����/��8G,��@���dU;�2^�+��E���>4� ��U��&�Կ�'���XlxVHYEB    b087    2540=X�Q�#F��C�&��vn�ڡ�R�{]�a�z����G�e�DS�R�m�V�J�����Rm���s�(��iaWf�f�y�"ITN �`�#In���,MO�cE�(5x����[87v�O��<q�!�K���'&��� �o�Q�$la��vyya�)�Y�m����aml��9�0d�
jg؉.�y�?�X�|�C+��!Y%�AS�D#]3qs��?��Ȫ���U���#�|�6z٧x�$���U%>O���!�l[�5�{>�k�p�5H�7�1�n�?�{��+;C�ʰJ!a�i���$KBM�H�&Z|��y����޻3�o�b>�R@�k���u8���l�mS}�˭tE���<�F�ƭ���cG�֦@���S�)W�n�j�Q��Aqr0��ճ(�
�ok�I��wHt������I]Z�%���"�I$� A0�8����ߕ��[����J���4MTBr�1�ϱg�p�r�( ~ÔX��d..ʩt��b���b�L[�	=#Zɻ&M�VÓ��`E�1��"���
�����c�4/��%�ξ]�]����G��Ϧ$b}�f}Myf
[�m.�E���k�a}�`[x�,��c�!y v*�G@�z���B�鋵�ި���q����R�����uV�e.���I `���I,@�D�t<w /���?��*d6@&�Т��
�}����ۺ�s`�i A"�D0 �16�l��S��b
V��,�)V��	˅��_��W���3�g�u���eu�6a"�<�i`���Q��]񀖳��j�1��2��`�]^�+[
����8p2CM�S���+���������3��?[��I�+K@��A�������Ϸ^�{ t���60^b@4� ��t�/US�X�HJ]-`�kW�P�_:�C����>}���~9��D�*�p�/䢧_�����p�=�X�e��)�$�����y�����M�����ؼ�C�Ec���8����ws\�s����p�!�JɊl�R��)�Yf�
%@+�6"����p�{��7޻ f�� _XD5i����U%�y{[�s�>�C;�������88#!�(��,[.�[��z�8���J(*����ݼ��ɭ��|fgK ��������y#�]ԅ�`{/-���欣�R����^�|N'z9�������`(����%�θ�	.vģ�k?�o�2���4j�\F���|�^�:bg�O>�$��/XC��Gy��`��7�U���i��_��js&8��|=� ����DAMO�[���U���i]��Y����X�I����ٟ-��m�̪��!�L��49��[{�#�����F$����Y+Xԭ�(0�I*��2a�1�j�>D��>���&cW���y�󅩸�ƅ�q�^h�r�U.u-J_�����3#���]��W����<
��P!�e,һ ŷI)7?�$v"�$��CAIh��H;JWSJ�x\T#�gB���� >����� ��B9y����� ���Y��D7�xÆ�AiH���o���e�� e�q�=�n kY����K���;�34*��X��)��>#��Mb�_ :��Kx�#>{�����͵ER����nA���,(
�f���Sch{�A�çU9~#�3��� �+|���s]�wE��� ��L�`L�H!pe��(p�%B��Jf>���E.Z�K�2��yH�^o"�,����
*�o�Es����r4󏞿�*An����a��@��.��?�7�w��b���Ee���q�"�Y�M�i�sbZ�բ�~k�S!(�F,Z2E;���"N�c�?/�!$��Й3h����f�#I��+N~��ȳ6��Mz�j��v�Y ��W���K��R���|���Fi��L��hkF:�n���Vn���t��u�t\׸��%y��,�5W�Fm���͏3 �^]�3[�wC�e�- �e����ڮa/@?�/�X�d�	̲�0�D�kPbO�Y��58�jg�ʕ�f��e/Q�|`! �ԩ���]K���|�	��Nq�2Hp|Qo�f@s(���@�ɏ�����F�CѰ#R�*{�Xfn���>ą������AB�g�%��}N��A�??͗]��kM��ƕ�L�نt����(��q�ٞ-K=B�ͤu4�$��S6�����lV���i���a�Z<B�ul����ā�뾥zT��_��3
��@�NԎE7?��q;�_n�%�{/�}��k��\��`��P�o��a*�\�	��εW�a�=���.���-!@�����P�WxtO��?i������C�k�j�M.E,.�����mE����%z��BK�>[�Y�WwH_g~���0��wg�1���=�-�k���U̩�p�����%�ɝ��6����.����q��UAz>+�f'
L��5��!���*�i���F���2~}�� �v�#��mC:ҕ;��ܜ�5���������
�ʢ�&�b�*����.тn���QXأ��q쨂����*B|�7l|���P�h &�q�5W����R+6��x����6��X��d���OlH$�+ lp���j���A�*�"sM�F�<H��H�f��l�/�%�(������#���e�L��l�Yu�7i�l ���|�I:k]F��>L���JT�w�7� ��=��$H{]�h\ۧ��\�@�wۜ������Dj+��Z�"�WT�Wr�y!�[WpV����ZW�Q�/��W��|8��V�)����U��.m��F����N)�L����m��eMy�����#I�b���(iK�*Y���??�!�)K�5lYL�Y���0����cE:a�Ҵ�"��-���������vq��g�2� n��-Z�:��kw�� 7n�� 7�h�@��J�&E5��U_Gn*�j�ԇ}�|h�E�����y!q˿�I ��?EW5D��:T�n�a�v�:+�Y�΋���~Y�y"U�E���JvӖ��w�J	@���l��!�|^H������_�q�c*�P�T9<C�ϨAV�����R�<�gˎ�%��H��$C|���o��;y��5�k#%��9��ҕZ*p3�5C�������B؟#�^���u�^�kRi��*QkP̃%�=�1[{��1?��;�+����N��x[�s��=M+�e�@�-�r�z�>.���qKd�� �t�v-��f��ܵ%",��>�~6�ƴ�UA���C��S���	v���+�b;��
�����e�~.��U����.{! ���B�;L(�����97Q�c�>�	f0v������ o@9k�#�'��#u��!b*��ΜT�Vҕ�ߌ;�ʿ=��p��	b�Ӈ'����!MB��h>\ؠ�tD:��ݣ���8���*TA�y��Aȣ�t�A�c��]�:=�p\s���-�����i6���>�brw�����F���Z��2ܱ4�՜	#����(s������-���\��0.i}�^
TI��a�_؝�����gڨ�w1m����k�Y�v����"��\s޿����k>��FnT{�u�6�j�IbnF�E"�F8����Lx ���W&��S�]��q�"��������ig�����P�}���m>=�:�)w������NNA�ȧvzc��P���w��d4�Ls7p�D\��7���qK��h�ݰ���e�&j�{�H:�O�J�a�����$k:����B��8!�N����N��gB����-5v娠�C�K����B-�"��	'0Q����1���C�Y�R�lY�iu �xDެ��;��O*.z�)��f#�%���`m]�U�.�㩈��W^�,
Ƥ;����U`]KZ]7��z9��z[�P5
�.
*~֟h�����RQ�k^CI����L��o?���b�Y�Z�7�n�J��&d�Զ��D���Ȱ�8J)IO���%E]�{��4e�O�Ƽ@��+*L7��M�7U�BH�ZY��%�_���$�b�?%���:>"3R�7/LH�Y��Xt�������}[-d8;B��һzf�6�㺽�D5��m�er��%�ad�x�M�3<J��<0�|rEZ��١�ͼQ!S�bx���y�D��9�*�:9ꂌ��j�WY;͘��z�!�{ZUwv:qp��!P�K.�+P�i�pkU_D0�3�E'h��2���'vp͵CNVʩ򑦖7�qqp&.ZqlPR`�W�|~oD�l��S׺	����D,��b�lo~e�
᭘���cˇ}�C-���D� ߯��ɦ���5���o'�����#�T��7����da����E��}f/��ր4a<��h��]�B�(��k�u��G k�:j6ڐ�z[Tˏ�=�c/c2YX���估c:�҈i�r'e'���>UU�/�.[��cN�p�s��z�����uG���A�A)Ҍ��ᰔ����\V��*�j��~������vg�lh��U��|��a�yMX��<B�����mrm-__��AwQ4UƛȐC��^�J{Þr���2�qЛ�eF�Y�����zV�� $ �0�E��j��ypz�Ic��5�UxbXY0v4F�E3�$/���y�$f8�tm�J
�݊����[�4<�M@�� Hi�s8=c�Z�1�SW���3�mRm9���^=
	h�ǇYi]J!���Kd�^p����!f���:`w��y��}�8$8��.��&3����?��L#-1OQ�"���3��#t/�L(ܻW�@ -�v\��P~Zz��Ln����γ)w#u�{ �LAF�pRZ&�,���k�,E�6��DJ�qI���;�ً�%�w�(�����Հ7Oy�HE���� �|P��W������ud��k�̝��u����S���	����TR�V���O=�r|A�r�/�)�3@2��ǺW����"���}'�p �|n���~H!���nw���@�Kʺ�a�?Q���~�6�?70�$֊v�P�	�[7"�v� �TӳXg�6����F峵p'�]]٤6�ܚ�;V�w("R��|���:�v0\���^a�(�ڕ#��*���� � yyy��F�']�0b�N����D_�K�׻��'�A3�u�`k�@���X�֛��Lk|f�ݓ�7�DdH�O����t�0Z�^[����V��702��U�<oL�BM��h}cu�Վ�p¬w�OIJ4��VC%S��2�ц=#�޺�*���-��b�Nm�ȬשzW����2
v���_S%���)�t�E��sy	%��8�M��orJ2<̚*��Q�B��d���ti�p�+����f���A�?�}�œ���R(�1a�K�#��%Zo�DRq�tÔ�����d]n��i��2�z�4A��K� ,�'�dT4;�	5Gn��r�T��D4ܔ'I���Y�i�Ga�b(�p�f�ңM
��1l�že^`�)��-<�fL�LJ9���.	�R�ZW��D'H	�t�����=�)1j!<�-L����(�;j���O�.0�3������9nW��\-�?����	j�י1�2Rm�2z@ׂ�r
$k �E��˫B<By��qe�Fk&u���H2��2a�H;���I���m_J�sO���G�(LU6�$�b�%�t����x�v}����*��@�D�f��W�g�����E�׿��hv[���F�T�%_����-c�V��p�k/&������X��7�kc�V�a���Ѳ�MFDwG�Adp{T�fQ�s��]��hdl)��:�I��vx9����#��fV�o][x��K��X���j�� ��,�����I=�,mCuN%ِ��r�f&�UY�����q>i5�3n��!�+���T��]�&��� L�3P}���H����O�3 o�C�s"�a�O�|uM�H�ͩ�n�:�L��2�d��\'�ۜ8�ӊ�(|r���1)=q⡝B�4i<7<�DuX�P��e�p�=@��;��ؙ��ղ����&���������,�q�/met%�t8>>kY?������kQ4q�q���f:���a�V݂����ax�կtF��hg�\��y�J�DE?�l}�#tD� eB�]��a�r��)���?����(�3}�-��-��Y"�������pt��װ��i�Dث���
�" &ͮNX��\j@~�F^K)���2�J�8����
�h�;���4�(Wy�-t/�ܪcp��ݐU��t��� ���؜����igo��D?&r��fQ�y�[�BC�ZPW�}���ӰC�ms�AL��YB��Jc�Vf{$�]}�Xc�
%�O��v`3E��$$�jE�_��:,P;���f�m��'E0�y�5�|��?���de4�`d�l��Ut$�]r"�ѕ����cMw�t@�-H�RwW�[��Ծ�`-�s`ط��"�����M9���m��(<wMk�#��~Db�&��,͞��-h��^n�I�4�]���/������nv�z�/�_��'yĶ65rg�g���|@�,�e1�����ӨU�P�B&��H^����\�A[��9"O0X���$�x F0醇x���g,�=�y��O�ߺ�O�ƹW���s2��:��~,b�b�켙SIi�0�S�q���Bq{�3��$���k ۄ)�Cdtu����!�8���.Di���%0�17m̳��ڤQX�؜����E��a��|B"!�¶y��� Z����F���"WMB�7�i�ZAg�����i�Й���P↥t��j5���d6� s���B��d
z��w��z�.����r�k�(��jiIߺ�͑��BX�s�����ø�e����M���y��J�U�[�Í�@x�7x�k���C�:܊�
��2����X���Ϣ@> �6;�uIi�ؚ97e�����򉃢�+a,�����5�q�͡w^��~�5�����������K<�/0�K�Xmyc�e&e�)Wҥa����e��Î���xc<��N	j��L#P0[��䊇'\��42��$��)*zg��m3m�w��%kn�5��R�����+�K��i����rL��Z��8�L��R߾�kNڦ>󬆵����wM�;yK�O�M9���d��3����ۜ�&D���jnӂ�sy���wލ�v�V�
����M���-��oc3J�C�������(���!�Z;�?d�4Kڔ�
��U
�I�.��*ڲ�te+�2Uy���>
��0l���?� �>���2����VқE���+�¥�?� nCp�F�X���|�!��u�������r�"k�$���T �@�Ec
�����#��ds�V%��P�EP�:l�$7��oy�~�߮�,f��e"���d$U!@�;�vR��,o�qX�L��w*X���W��M�jR���m�]��ZB�B=s�H4����0��T_��w��A}�{}�_���i|�����{����XR<��C�;/����g����������vpGX�z����[*bW���9����P�ض;4,b���u�br�@Jgyu,@�%�.�O�j��~KAc���+p7�f���,�E�o��z;���w�Py��M��3�8�-��(��p{���2�j?��l�Z�	�mX��)��� ���2�
�A�m�����u�m���7/�k�i݀��`��W�T��,ƍ��P��y��?-����k�R]�h-�Ҽ�I��'*DF��G�a�0�ML�q�c�_��1O�D��ܥ������{/iƜi�ݪi�)�&�|��2�T�6��&�m���K���.�v΃�|��j��n����a��?����M�����Uiy��������a�mo;�{WȚ�����/i}os�o0q\S%�Pm�+������6��}�-L�c@li;[�ݝnD(�"�Otc�w����h%���5����Z���ɤ��i*r��ߞ<�wY�a����f<�W�?���xe��ŌR� ��X�tb7����\��#Z�?�d�K�f���#���SJ'~�z%�ϥ�H��f׋Ġ����wa�;7���NZ;�@�կ�d��+��Z$!�Y�{$g.ɯ��v�Or�!�FiF�"c{��*�5����Qs/y#pU�2-
Hn+?�	?��y�ֿ0�U��3�P2b��*s�l�|�3���s�@�#H��J/Q}�&�?�:G5ֵ����v�?�Q��h���M�&�X0�E@L	�a���g�%$Ʀ������Ֆ��2��6�9��)�>��k(���:��z�L�@��b�V�b+A�Z���_G`�~>8�]yHc�|������HZZ�Ӳ��n�<ؐd�4N
����=��������v�h�a�n�l�ߚs5���P�JL噛�ə>��T���ä���w�����.)η��@'��fR�M�&ʣ�'���J	�X�����Mh��q�+���c(q8<d���~���o�pCxUE�B�]���m&�X���	뒾Z�H�`��#l��#�"�Ap�u%�p�<׶ɺ�':�b��xh����w�Z��7j0����{�2jrFhK���=�y��+zD������	�	h���ZR](_B�����E��h�ߞ*� �:�*��GS��]ܪ�"h�Zv_	��Y�k�o3���*A�,�Z��yWęWRQ��Sԝ}G��Fޖ!ڈ8tgyav�.��qN�gƭ�#h��2R�� ��(�6���p}g��5œ��$�"YMuw�	cgǰ�ո4���9�=O�
���^�|j!� L�a�X��} 9Z��o�M��-��t�*���M_"�5�<�.�q$A����Y6i2��`�}7�) @_�adǩ<c�VAK8��3���佂T�p�$�T���faE�J��p���p�I5�ߦ�񘈼`�>,�����閡����C+�����W�2�nm��D��<��c��e؈W!�yum�����05��v�kI^�P��2���HO���RG����J����d�E�,r{���Ѳ�s[����_�(|<;ԓ9Yzn�����K+Wt�KZß����ѧ=�m�/���DҖE��7��@�ljl�z��[����I1���𙞧_\�.�Y��Il�k�7Q��3݆q�����	�kk��ړ_�wq��͌=���Z��%�'6R��0��dUm=	�I���y^���X���^��jk���^N؞X��8s�E6�����P�9k���ˀf~�)�T��8�hR�P`�a\����H���6�L��I(�fH��H����R<,}�7��%�Ԗ���e.�� "��v5K�y<ߟ��J��?��ёsN��{� f��n�Q}�p��Q��ʠ�g*4��