XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8���V�J���RĞnȢ��|����Q�+M�cѨ1�p���B�[�sYf6h��MB�浌<�RV�o�N�Y�'\�L-��z�	M���`4�kpw����8�P��&A����<N��D��B��z�`M$�Y��j8sr�-��g c����]S>��� #t%�����'w��2'��1�HN�&��dE0����;mp��^w+]B M.�O�d��k���ǔB�%1����Q�DB�;�Rn����!�˸ks�|�^3	_��p|TY�%Zj���͍H���?"�|ܕvU�sFg	z��47����Y�d{�.V���h*a�#M��0�����kZ����M<�
j�x�Vcj��Y-Dp��|-�c�k� �s� gy{I��-U��X��}X&.�@�L�kL��F��v>�����@R�񵬙WZ�">�w?����ɬ�2O_��3ޚ��#�I��/�����0g�jKX���"����|ى�\Z(��$�4�xN���ZHta��N,]6�A�H��߬p^HV��؛�P�
7���5o�"w��~���o����!݊��7�rtf�Ty����g/����}IW��-��C{��}�v������Fx�\�5`��`�����M7�0l����%�n�%`�'ѳ�8�X��T{�גR�W���P�9�u�1jV���ōPZ��_~\7?�'�����kY�&��'P%.����q��o��ŉE�!b�D���[a�*B�#�d�~$�kl����j�N���"�����XlxVHYEB     e07     680G5����`��<軤��r��C
��V
�۵�����/07��Fݪ�����G[M�ҵo'�RU�S��ѺS�i�q����l��c.:�v����>�K�("p�,:׀CCU�q���t%���Ӏ�f8FF-U{+/v��c���CH����?��� �a����fq��υ�ۆ̬
[� u^xd~�s�C�y����N������]�Kh�3lo�=�L�� ��b���ҍ�;qǗ\�ޣ/<VӒЮ��m�^{Nc��җ:.1�ȃ�����C�Q^q�T���R!��0�V���`s(9U�Pұh��/�{�2�~����H��l�c?�t�O���ׅE��[��h�miי���UScȓ�o um��4���X��{�14� ���x�i�Y��/�S+y����24ogݤ���)�p��Q,��H��F`�;�ת,PkZޥ�[�r�lN����'���9M� 	"�iN�3����#������+� (a<�񂃅;�^_��b!��I�!H�QL��	�����k)~�L��]F�"�*p�;�D��$��� �DJ�0nk��q�/�a�V�x������<6��	��������
RbRϭ�j:�A6�?D�eҤ@G�\(��w�L��]��x�1S �6�� ��>Q4W�IL��dݭW��z{��0��Hle&� ̨������&ȼ~��I�y���]so��p�\;O?���^��e&��o����H��b���$VşJ�v�$'��]K8U��Y(�{0fe�'�?OG�Dh|��Ò�z}I��b��h�$��@���ɯ���~�J��ӕ�����V�m�g�3��|����EF`��e���ǔ�)>�<L)F�:E��`!�� �B5���N�՜�_�K�b��zV�ڪ�q�ಹ��<����_�*}�J_v�`x��.ɡ�Wx��6�G:�D�(cN�����p��/�`�<�76��h����²���\�C`��	M�H��&W釭�D�U:vΒ��F�+�MIed�����!Zx�4���񪁏t^��Z����� ǥ���.�Q��'��(�E�z�UƐ}HWZW�<i�ex�ᵱdxYk��U��1J�/�?�LY�jA���f`�FV�1;"����x��:�9���y���5�E��Ԅģ,�U�~Ev�T�n^6p�[�Ur�\T��g��a��]|�#V ��tb,A}����� ���r�z滒��3�f��N���-��h��@��pF�m�x�ߣ���Mknt�~۠Ix���Á¦����u}1����u��E�()���;y�^L@%~�'����e�3�t�ڸsyt`~�;��ؙ,��z'e�vй�ݴ�!bx�"�`DB9��sW�B��cLG�l�"~�翘�stΰ8,���So�����H��/O�-3���e*P��X���P�(�'@�O�����}�����C�P���8����1�w�<��2S�d)�%!|�P/�:�}�n6폞]`�{/����wш�C̅�O�6���?��%�{��p�Z�c<�ݐ�!A��X@�e�y_��W@D�k��rʨo�\FN$�h��d4J��B�3�A,���F�01���Sw���g�a5�=��'!��`ބ�