XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����=���LT���N��p�
��8�FX���
�iSbȘJ|PxU���{��g��e ֞���N���'�g��BH������:̾��EkW���H�Jw�y��]$Ƒcl��d#��-�Y��@��z#K�yT/���:i�[��̙�*��d�HWq�5-8���8�.g\hdq�v�a��U��]�U�뾰�t|�J��;�tW[���y���9qCbUG�Pג�({���qy������*��T-H6.���a����כ��d{�OB��S��9���f�oT���a�m������ⳅ8{�6���a�I{�� =�LF����SxG�@d'Y�k*�����s�9|
yBi�ub�^��b���zw�D�^bD?B^�H[�d�����낗�q	iW聊�ci����Z����ϹNO�7$aG�e:�$Û����3Z��аs��+*�� �K֣=���yKKڕ��)Ea1�-ExŰ�1p��y��S� �������z.�{J������M�Jk�(C���$]�s&Nr�\;N�z9L��s������[VS@�_��*t�χ�>�@gR4a��M���q
k,+J6�j܅�~/]¤���Lj��k� �/~!d�!\���1q�=t��t���5�bt3J�[�O����fH쑌Pɺ�"�C�m]������-0}�X���;�o�HBA�'<&���ʏ`Ħ���e)|����d�i|��<ց$����IǙ����Jɰ���=�W?�1Ѻ�pXlxVHYEB    9fc7    1fd0p`V1�
L���%G{�*!�B�UCH��ո|�C�L��jY��:�̀T�>��vS(�D�^�"�R���a����h=�H�*%������
D�jG�iA�<�c/��*�� ���F��Ę��8_���n����|tNI;������~A}eƻ���KA6g-��B��B��k����}~&����=r��)Q�y|�/w�2��f	�\]�t�L׀2T�i*�����mC��(��C�.�_�8��w.>�n����舏O�P!)���P� ��&�*�����Z�+Ҫf+�:V�0NMD��\=�>�9�^Q�;-Hws4������u���)M�T����
�+�(y�
�Id�LE�W�{o=Qa�\q������1��F��9*#����Ky^0 .(����)�I̩���� 9���
jˬ:�1��ɺ�=a��UG���Z>N�"�?yu��X�c�f�$ u�y)%�V�9�r�J��Aξ��v12���M������; 2��
լI�V��k������h��S�n�r:���� W��o��}���|�0��}��yxc*�U����h���W��lpX4����".��+�']�{����as�!��#�u�.�:��L>�(��Xߑ��z�&(�=D����)v�J'�.�����2�{�jI~��Eh�2��x�L�ia�:�X���\��+���8�*�,% ��;�o�����"��j�Ď����89IkdҤN�E�NMGP���V��p�1Uܓ?u4����(�mţ�20Jv�(�r{��m��Ԁim�{|��s��5m�r�&Ÿ����=/�&��B��� �O����Y��H1�"t#�1��?]f۟�r��n�Qbo�xC;A�1{,��2w{��I���p��>�@���FQ��څ���#+�"+�G髄)����k��������gA��L�z�����n���R���`q��~F����~�P�过h��o�ݙ�k�]�XJç9i7��07�F�{Tl���U�_"���nw����ۍA&���uo�&��j�曞|(��zI��eN�`���ޥ~p۹��&{ւ�PD8D܆(���������=	����+��eO�+G�5�AA˧s��M5�����ҕ&�p5
��.$R�������ޡp��TJ/�gG0���D�0�2~���l��y�J�=c�34��}kR�����sj���G�{{<M�K�>�,1�a�/+H�h��7�;�K�7\��8��Q�H}��V�k�ŉ^@u�a3�����gU"*�H�(p�m�Ƒ��?��������"���uf��k$��^߬h��Hv��nO	Qt�#�m;&�4�n~A��$�cQ�.����iA���Ƿ���5+7��X�7�w ��hW�ʉR�G}($d�Ǫ��K���9^�Q��h�w-�T�8�r�\z����6� sUA�']¯�h/�>m4� � �$�N(R���+s7D��D�L��'Ees�ň�i"n����z�ħ��f���Z��4�)���~4��۶��v��W��CHH��i*����E����"_c���e��G7�nL�q�`��a��C��x���rF9�S/��:kߜ(�0\Jx�i���P�rh(
;�;�ܫ��������OՀ�ؒ��$4��n�݄�+������-}����$�zp4�޶v��7d丂`�1�9]���T��0� �$G�U)�]�{ UAW!��{v��?�Yy�"j+!)J��J�'����k��P�K�����C��'"[
�3�<h|��8����ٮ���m;�s�&z���2j�����1�� ��[÷���2ƈ!o�Ǩ��=�T-h��o�u���>�௕��
����[��F|b�t��<t_���|j�~ ��V�L�"�|�6L߳��)d+)>V�d�9�������`��y�n֘\Eg�2����X��٭�J�K�8�C��
�(S뉭��6��cA�]ġJK����%;	fs�}G�ak޻�\�|�p��S�δ��tg��S��d�eRٲ��/MM+r�������4�D�{m~K��2n@L�Cӳ0��I6"Ar�ԼZ̝�00�]�B���!pb���F7��?݃B��d�Z_�	��P����v��^Z�C�FS�Y{��r�6x�F�|0��f�e�k ݋
�h�Q�|�F¼R
�;�<ouP���ҽ3��T��
3l�E��t,4 �m=]�e��8k5��D�Sk8�m��!`��}ǆBbK@ km@�rc�7�S���^�&�P�����/�Ա����)�#�Z���wU���3ӵ�Cج�7�ƹ�+p��o.bux�L�w�E�����u+>��$�����LLgK�EA0�zOty��nx��}���)�'Y_�����- W#&��tԏ�u�;W�<WNJ�;k,��r�eX>�
止]�%K�+�1� �`Ƀ�6#���v����I�6tkw��!�}�	/;���Q��� �BN�\*A?��}L�÷��i8~�W9%X��Y��M���BQ�<&�W��:(>g�����lD�H��O�QX"u��&�#�𚗱�O����[��ƫ���,��cǩ���^�Aߝv�Y�I�_[x�f�����9��"sS��[�Fx��Xi�>�����,�3����D������e�����_�����4�l�i���Љ����-+p	U"&���VaH�,�3�r"���6b�v���U�M�b;��Ǒh/�����%��$�o�&�/�y�����!�R̹h���P�&}-NE��j�$��<X�4�n3���$�=�P�ٞ�^ҕ��`)�����E쟟g��E�_m��,����$5��G��B�������ڿ[j�"x
pQ�U*�=E�N���1J�lbk�y�V���6{:LG�Z9��;�4Q]MΧ�G�lg���2��k��*�x:���O4��A����RdD�^R�AM�֜��m�-���4�����+ '�F����y�X�*��q�RM�d���E]��&�e��b��lH�@o��aT��芏���H�ås>�:6w6e���S,��m�GBM�|6��
~������@7^5#9��RҜ���
'�L�����f�s�i��/{�]Q#�JՇ��CE[k�*"|�E���
f&��*�V�I��n��� �E=�98Z�yl2�A�.S�x�m��moi��꘬���ŞA��F�Ϣ�xR�>�$c��(�rb�d���q��u�[���^�c:*ܶ���l�=|�
+�F���ƾ����*A�wll�η)��9�D8$��j���a�<�|KŲ��'�mKRړ$5�A����,�+�JaƼ�e�����G9'佂�>��Ryy�]����7�y�I��2���x y�,C@��<%�ˎqLj���
j&���k�H����ĸ���s�QuD]XU��w��<����/���3B/���)����'�~_ܹ�োx��T���/��#a6Z�����<J�����Of���y���+5]��"��c��W�o�z�⠤;��M{Z�'9�'�>)�C��?�������i�Q(�z�����J�vۼ�G�)I�},j'>,&�I� y&=�d+�ܛ���x���ph�?�=fq.(�����Jq���ة��By�1OG
�����B�n�����ԷO�M)#�Y�Xi�����!ι�����#n�~|+�-�͌&%aퟳs�Xy�O�'pb��TS��m��x��w!�]�����󝮨�AB�b�>�DM���آ.����/^��h�	��N%��1��fB�}�²�pO���orii���D#U�]�߃jɋzX4A])�z�VqUB$2�(e�z]w���+�|�J!�!7�Q㒔0G=�[�0�̣�k6x(������E��CӦb�u�n`�-ۀ�c�؛	NE�B��HI�a,G�[4ӤK1�U����i��$�hgI�.���Ȑ��h���)�=����`�$�U�(R��U��?��;�&����APm�2a�Y*�92��U�s���9Ԅ��a�,��μ������K*����`e�~�6(�8K���dQ�E�=�Z7O�y(��¼��O
3I�xe+���Fd��`nt&��x��,���hf�p~T������b�q0��A�k�;�r��$-!�eZ�V�t�2-M��`��B<S �Le0y�$C�{�p�xT;���+��9y��Ki,��`g���/�%�#<m�dTf����;gT��c�b�f��PG�[8l8���/�R��t(L���=���K�:��$���D�5�}�d�yS���
��L�֝Eŏi�3�޽U(ӥ�����X4U�ʌ�+ �G�ט1����`̟������ǃ=��1 �����-u���m?;4
�������L�h�Z��x�J�o��=[���=E����J���*v�AY: �1���Tq���q�`D��E� y��|����8�������0�#��������=����I]|I�3���S�����}Ⳑ�%� ^�%��r�P�Q+Fh�����	�(���7`5����f��h�6�UY߹C	������(�I�A��p����縉S��F�eב]�H���R�mԠ��w�BEW�Jg� �S,�{]�sUrZF�J�?��T-K��Uڲe ���,�����B�� ���o�24���n����nc�zW z�p��ޜ�4<�����������w��q-%{�@Q���G��kO��Yn��zR�1�,���ydj�6���wF'J���'���D��+tި�%RY9�jm�����(s�9n���N�8;	��T���"�V�����G�]y����S��I���I����u�N����o��/�aw����.\��I�~Y�A�p�7 ��?ʔ��
���|J3os���� D��lQ����@�-kF�/�]�\��Loۖ�*���S��ګx'����-��ؘ�.F��+]� �hxR�q�C��b���rD�����$��I��cnTck�㶪��a��:�Š3��I�tu���`��oъ�O�=^��	�(0�AnV^�~w!�E�3c)�т�wH��`��%�pp��\�@�ru�P~O18v/
�Y�$f��a�ټ]+(F�r3�<C��'�g5���|���*��7Hr.S��p䚳��4O�E�L�m��.��d�~J��A�v�!���{Z�����uf��Q�,��L�a�ا�O��:ɐ���jd��"W�(�M&��YR-���g� 4=�]�ұ����uoL��2�p�:|[������0'�U�IC�ĽB��|�̗|/@����,�ZV7z�����e觗��~[;N�Ou��VhW0�Wd�Cެ��y�,0Ax�p��p��CVR�.�E!h:�ě���͒�~;��	D2����8��0�nʆa2�k��%���ļ"�ݿ�y��)(������{������?f|�:QO��sӢg�y`,E�w��'P��Y�a�%}����oQ1<�'�}o�8�5E��0���#�Z�G�#���H[��#"��F&К+q��_���5^_}q�J�;��
��RQ�KtX%��[�����յl�*c����{�hO�V�y|�Z�ĺ��po�����b�mj���u���yc¦
'-\a�C���0Q"C�2�͋� ���LW4�?m��P
�Lחጔ�����V�B���8v��f�����S!k�!� �9#��h&/��^@�c�ƕoO�X�6;(]����.ɨ+?��Qj�Z�ì�osK�Ʀ��23�Lu �a9 �/����5����F*ά&�Jbޤ���2�(���x�B�V���L��xky�a�Q$%�͏��|���j���w��|rL&�
���XѮc��<��YB��I(&���B�n�hp�J�T�y�rʮp���������ª�c�s߁N*l�f UG	Xk���z�Zd�xe���>�VJ�/?�����'p��.h��߇��-��IV!Q;;wf��j�<p2���h49�b�]��39,o���$���� ��M�Z;�b�B��-���A�b!S���s�:���1�*<����Q��>��c��}�G�;�v�cfӠx����Il�'h�k�z��Ț�ͣ�~5��L�|��6nR���|��m��FV�q�%A�;S��r�uHaڼe��;�*��-zOd1f.��=��nØ�>Srz�x
�0�ٹR*��נ�H8Ce�cs�["�n6)��	3X�8��!Y-������NQ�ߛ���u��#�<3���p,�{S�@Z-��}/J�
$�p���N
m^�Ƭy��y��Y~�ON�Cn�9i�o���Ŋ��{�I�R�5@��������u��,�8)��vr����B�����`V�p�]�%x��7>!���	IT���>����|{x�}�U:ԃq���Q���ȈKn����g��ݤɽne'm��=Hһ��>�.
*I#���s1��k�{�����=j����qm��!���Y�@�s�ͩÏ �7��$߁Msr�� �r��<��3�ڰ��"�T�9�*�J�.N��DG�"��vk��ٕ�T���{[<ӿ��S��� ;�<�<��&ŋ���mꂔ�3`	4�M���Q\��b��3i9C��=��[��M��z��Xq�O呈9����E���8J�7O�f�=	��_A���T�3+��M;u�H�>`#L�G����*��@n6�Y\3��|���Ie����2��>�Gu�hyv��W��D�ӝ]8�{�vQr���4G��si1Tj���:����GԠ��;`��!�Fh���)�r�5	��_���:����K���F��j�����<����9�>�v���O�i��J}�d��v�ԥkcpG0H�N4�}T	��`����#�A���;�8���=�d�u���{�Q�o�T����̪,����5d�Y�ul&lL�]BwhL�#	�X���w�����ͷ�bTE]���(G�M���~��f�i��z�賄��m�}���F��CO�+Zn�V�3�7�6T�Xwu&4�'9`�}%+O��b�L�J���:xLA�k�/r/Q�|���g���V�Xw�q/���!���n�]����[��1���J
r�H�<��R>F��䩍#`E�pt����Èx�Ι�N\�9��5bF�C�0���L��
��ei��S����� �eA�vO��r�aH-7\�⾖@ ZcW�^Q���DהIg�����bVrtY(z�tv��eO
�����^]��R?��+>"�8������ku��ѧ%�Av����+�V��:jT?N�{]3��IT�&{J�~\�^ޥ�C(#��لKꘂ����ԜԀ䫷�0����#���1�l�>M�e�����	˜{4;�,���8�k+�crg��4P0@��.'-�3�l�����~fd�_nl������@|5�Ё�ð3#)ژ��A; ��L�[2���P&�N�R���d�m�c9m�Yjn��!���9K����e�_��c�q�^S�O�J#�I�n?�޸R��y8��mS_��cL�Y(����[b�y3����i�m�,�^�ihh�p�_?=�~d+��HP��J��)٨<�1Ġ�M�Om���H�H��KTY��B�&�� ��z���3���^� �*T۳ٵQo8?�OWs)j6S.���}�/?�%�~hn�s��k/����B��u��l)�ꪝM�9O��)����j�|�b�}�2�s����J:ް����~����w����<�y9��=���%SP����E�WL�U�[�U���Y��ً�om���
�(q^�rE�{�a��#��w�H�J��1���aY��׶�A������M0B]gi�!�9oY3��غ$�Zf��ͤ1ћ���JK�.0J�I�n�)���ގ!D ��kzA��+��;f�o���4���M� In~��