XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��q,�����G觖΂S���Huo�-!�j6�{�f�u�d3q?��^�%Zd��|��Q� d�ϐo���4�h��8n]+�؋%���?h�o�jqi�f74�/G�� �6O������,T�o�l�I���Vk��L����>i�Zs��|"�Ό�ܱ�c�'$!=S�
o���:w��8	J�T@@`4FT�ѯ0C�q�y�}S�ͣ<�w�� ��d��	����S'��f^��e�ָ�9j�%���p�V�}p�t]o�#_���ݴ�V��K��&W��w�^�?"Ƭ���S;�Id.�vw�d�y�o����
����r��T�ƚI����3�|t�b$Us��x��W���e6�
�34*JE宦iIX�(d{pb�����z�M��%��01nh��*��l�9K��,۲9��tazC�{�*MC�Ւ�?n���d�e�x'���eEm1�oH������f~R������ſ���0�����C��cB� 2�o��v�&m�6Y���F��L�Y$(ʷy�{���)��O�t�4h����0�>��Q�'�>��;`dPP�qp�z�7�������m6f��U��'�&�N�q�a���b��tG7t�o�}eZ|�%�;�_����PsU�S��/��ӊ�n^+���g��lcw�����|LHP����ׁ��w�!ܐ���9�_����c��B���m�յ5�Fl-�s�|�GPF�SaS$�7��rMnd�ck���y�ùXlxVHYEB    3d43    1030eGŦ۟v��$]W}2�h����)K34};1 wPR�����K�_B�ʧM/�v��X�N���K�;G����yx$����,��4m��T���.���IZ���O���!ll{�i��0i��15u
l��D�DƷ����
�:a��/�/�cf��-��̴�#�DLs��B
G=8v�U:d�K�1w�&� �j�����%����&�M�N�:��(o����f�b�0�d���p��͂��릣�n��ʷ~�(����@ʝ��
܍H������$VFA({B-Zr\�Z%�����As����f�<=�b��Z�67�^��)�X�<��s�<ߥ7u_c��!�����{k���R���K7��UW��~,�T<�k�I�wX5�.a��FP?gT��kOз�F��s����Œ�o���o(`���pL�k������^E� ��t�s*-D���q�� �ڿ!���xYG��Ei��R�8\uH��t.�R�mɊV64�g+T~��x�|�ք�����b�¶}�i|!�a!<�?2F���B�|߻����';�Y`�ŨOtЎ�GYz�elȫ��<�B?��;�V(d��/ac��h3����
�ƯA�\ꞁ�LI��<(�m�吘��A���|��f�Lܥ�"4��'>�Tf�I�����沅F$R�{ӈR"�sw<#C�
����Y&��_"_���\�;38��ן��~Y杧�����3}�{7��Z�H|V�5_�a���3�����"��022�@�sg��	V|��f�I9s���.��wPs������%Z=�b��|g'��k ��hR]:�t��k�$�L]���+���f�&66�ۂ$�
	�<���Y�y�9�w�g/U�G�{j	P0��.�odʉqN2��Ku 4N���;.�d_ �B2� ������`;.
Q��n62h������o n�fuW��L�ߖ����ς�b��ug��'g?�ŋyn��AC'GH�}Dx=5�<.6O�?���.����`�-w�u���A�T�� xZf��k�2�\V�O�,�5�^Y-� �9��������V��4�2���
w��C��N|Z��R�0u��H�2��)��]�F�owx����i.b�#8L!&0x2�8��X�t]4_&?��H�qr�f��}�P<��.+�8yƽά�>���;芛��(H�#7G����;(�p0Qj-��O+Y9��	ȩ�����=�p��w���C������"m��Xd,yj&�i���~OEa�����~�[t^kWj����6ǻ��9l9�]����I�g�9D���DE��5];b����]�@3���k�kЃ�8���<S�ب��ˈd��������!q��x���"���1x�1�P�0`�/u3����e=V��0���ueI8JY�DqWp�U%�ax�1aȕ�Bә�g�1	f���(��J��O����z��["�����%��΅I�w�Q�udLB\�8w�5�0��^�0Us'ܧל��1j{�b�2~�QS����x�/�/�)�9���qm��x��Ǔ�`�����)�ػ�Yak;���t-$J,�G�d�\s)��0<Vw�r��aF�a�9��F�^�\�E��*���-��dY� ݚ�,�4�YSQ���5�k��y��	�^�R��?Ο�@n+7ס��V{�ϖ���k 4-�9�h��K԰(X:z�=N�M�����PȚ��r;	�!L�p�5�%a�����-�A����c^��q�P> ������R��>:*t�XJ(R����5I�e��O\��
nL������:��Q��m���٫~��u��@�x�c��eʥ����EAfv0ن���w� 0�]Rz؟a��1C7�n�Y���y�n
��V�� (c�sF�.PLiO��i�`	�MX�i���TNR\�<�9Љ���o���=3����J�ɛ�u�u+p��=N�e[S�^�W��A4I�>D��Χ�rS��ݦ��߼�W9Hf���j����L%�d�B���ź|L#&p3B�i\C��H+=�^��qy���£{Ֆan�f}��΃�7�ԟPK��=o���E��P�9���AT�킣��퍃7em�+�������;��	��G��@)���ױ�^����[F#�W�vʀ�������?�}P85)������^\,,��U��#��)�ׄ�I����MiE(=X�\c��o�t�������|���/�2B�z�n��T�����\�[b\���Mٞ?5	L?��Zxj��:�H"������L\Н���)���^9E�c�߄�{�]B	0����l�O��S��n�+�͝2����xL�ui6k�h��$LFB����{� ���Ĳ�4Vj�<��[�Ņם��^�*�a�E8p^�VFC[d�S4Dϱ�aA`�n��'�%Q��ig&2穽�
����x(����Ϡ���BF*54wZ�;�jJKg@-�0���*��}(�Ն�v�z��><������N������9T�N��[ȗ<F�O��t�5?JxA����S�K��E*�|j�F �d�n�+�=Dg�_�F�ê��-����fz�$�t�� O�-���T:'�b�y�пtm�ŋ��q�H,�}hK	ɀ�/�e�G��f˼���\�\�o���o�-�O �"� r��uůK6��P�@W3a)�ެG>˯&*ஜ��9�}���}����r$�y4Iն����<_qa~i�����p<a��v�R��.��S��5�����o�l�e�jĎ?CWpKD�H#�����N����s1u�'�9TcB}�(� \f[!�2{�G�D��_&�����)YN��ʁ�	)��L@;�����(�d=��?�`�0Q|ȧ{@�D68-Α��ơ�#3P��2����'U _��R�&�G�e`��3��֍{�'(�T���o���D�N3�6<����LD�!��4��modJ�o���3�7��i��e�ڍ��1��Ξ�d>��Ύ�����8�S�d�Y�hDF�a�Ϯ˄,#j���lߌ�6�.b�iH��.���Q��I��Sz(��}���h*����W�����B�	��	-C���n�%��ۂl��nI�<=,�����C̻����
������1&�es&��0�[�Ti���2�l'h�`�Go\�k�}=�J�R�B*�y�"�D�G%���Gp����M����[ˌO�y��E>;Jو5Q����2 q��v����5�vP�m�~G�ou�X�)�(�Jë�8O$<mu�����VKgu/
��I��q��!A�cA�Z3�P�Wۃ���6�	�z��?&�C�&�F�ȑw1	���D�Aܯ4XW/�:f�BV�P���9��_"zg�Uxq���"���Y�C�!K���Pu��e��Q"�Sc^�B�A�@b��SHh����Ȑq�Lz��ТX���j"�Mw�E#���N1��<�m�F6���S��59�/�1��FK�OQ��D>X��4~jX�a��go0b�j�6�>�m�L��ν$
�Qc�+�H�Uq�P��0t�6C�xQ�ng|pQ�t)<����(�Mqw�~��pU�XJk+.²�D,�,R����D]IfϞ�����$�2��.++�Ǔ�d��0z��f^�V|xK�-�O�`�t?��|nG����9b��<uuNV�@J�����^��둙+�1By���u�Yc�X�뽽��ܪׯ�@]QQ�jx[�I���t��l�"@@8s ����{��d�9_�yB�%�`�<���/��-����A-�k�c�U;���-湆��g	�p�vD��HFl���)�P�W�	Q�[#� {�������XFaX�>$�vO���3�Lx��v`X��Ӟ[��h+�����L�6�Q���t���64!��������|��Ԡo0H!bD��/D�G��;vT�N�ʖe�����>��n)'4�������n!w��H���x�:@�o�>���nrA�������/b�(5eg<�t��Gw$Ni
<<띇�E�%�7�]��c+�o#�