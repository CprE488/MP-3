XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������X�E�`hs���2�F1Fe^X��]E\�\R]/)�x6	80��Ŀ%�3z����N����1���?Ib��]��v����gJٳ�V�����j���Ȓ�2*Br	'�Sє�V��owy�{�c��N;�Ι�T`�]{+��	����xc.n~�Dw�ˢ�$��B��[3�B�(M���[ bd�+$�5e����xG���7��4�b�԰@����zs#�ZLD����A���2R��s0x��	�����i6����� �j!�R��ޜ$�$�c}g���yW��
2[�'���i]�X��^t�(�ќ D���92��Y~Fjz��S����g+�|E����ӏ��pvkA����>�Q4t&5�#�b��(����i=��m/�5f�^~ި����i�̦���	������s��|�uѸ*K�5�0�Pʄ��f�EXo ���j�c�#DZ>�e���ݥq��&�iU��A2#�����ܛ9��k_�%�zY~9~�юkB�&z:��9���#��;��:@��,����?e�^����6̬L�
Ľ����˻?-N�jߏ냁�L�Ru:��٬����r���[a0E�2��6��oF�c��D%�U�_d�ت��}����e��ʻW��}r�hC@�����l�3����U�#"�:���;(D�Y�թ�
�mnԫL�N͐�Ƌ��b6e�t�-�Q��oSҽH	��9�v�?�M`]�$�=��oXlxVHYEB    1853     810ѻ�	�oQ��is��f'P��PK[x~p���=�=h�z���P�8b2�/�2U��C���G׎�!	��%S1۱�`��~l��m�8M��A� D�$&Z�R��'��qq`���S@J/�]�7ἊD��S#���;�����`Zr#)Q�b\��0�6�x@b��p,�W��\�����8�F'S����/�W�fTj[c/��]���Hf���\�ݫ��h3��p=����36��q�\$4��\��Q�4T�($TΩ|^	wTi��%x6���ٴ�	�@j�����K"*Ҩ�%7�y� 6_�d�6ˀ��l������t�9�I��m��Cl��n��.TFL�D�����@L'H�rU9�= �6q�@�8��uzE8��;	`� �W�2	ܞ����vN��~����$QYE	k��;�B
J.g�O6zU����b}��
8H�#H�4�^��Ӊ3,r}���9
$�a�,J���)O�Rh�W)�0Gf��u�G�'�֎4��p��v�S$/�ڴ�Ȭ&��x�r��=oٿ/��g -��N+6;���H��N`*$�S�q�Ux�w6g�~��-�S�X���2�4^�}������<q�WԎ��K��*!Q� *�;�i���8�zu|8v�q��N�:���B��N�X��R�������(�A���vrM�V6� �Q���r|d!-�Z#�1����6�"����*T�Q+�]�r7Y�Eӱ�(�����S�$	$\�B]ɨ�$�Os�tw��w�ɋ���k^?3�f�Jn�č�����*��^�:F���Ptҡ�����0���4=�6�.k[D�	�+��򑽃C�R��BI���f�
l$<*<E:f�x��.ܳ���i�4��8k�k�D�)�]��i�A��dm���5_��i��4�3�=��l�����D9:��6[~K?&�J��6v� ��҇v1\���^7pD�L�?ԗ>��������(Y��t���j�8R����;��{�$��ڤj(��Vp[w���[Ho�C�-z�����
H8��Ͳ��d�
�PZ0�bzO�*g;m�F��X�-U��MU��j?�9�꼼�O��E�S���W�ގ��4TY^ ��j]إF�gX�}�b��^Y;����N�v�W���{�� ���0jR�qڷ��`����8��O8s�tд4��W��kx�K��Ӡهo�9��]�U���nf끙0N/'��x,dh���εu:Ųx�9X�A�}1��nI��0�H�	B���Mr�tn�&�O)��aОj��g���F�\-Ȓ?� Ɠ ٛb%�wc���Wv�'���4��e;|�r�J���beZ߼h�����ϒ�T�Q��PB�
5�q �٦h��&�I<�J^�F�ټ���A2��r�D$0����^�\N��W�Mz�k��?e���k�f���%��C�̭��s���/�`K�)�ÞBJ�+�H7���t=��
��×Wx�Aݪ��̳i/����r�=�������+8C`����'������..�,�I����b�Usv�60x��w]���|��^��(7�4r��=y}�ņm�����Ք�� >n^X�3����J�����D�����'���𬣠&�����St��������j��d�-�W���@����=h�9+#�ZOV+QW�B��[��`J�	p%�A����B1P�\K��x�y0�(*���>��+M���G��
��=��|�c r|�u\E��$��� `ⴡM?E:�6��~���"���S.8�D#�T�Mh��PuJ���?D(1�9�Aj{���)��̒��qn�+���-��B��1�#��z�T/q�k��P��_��'3U{�~�t�5�
N(k�W�B]=>1�
�iގas�d�>E\��DAb#�5�3���L�'g�Z1�cw���͏&fƊP���"� �9��<�bn�y]z�m����<}1�?՟tYvmޠu����� �Arp��X`6�Q�