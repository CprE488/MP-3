XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ҳ-��F��x����f��/�2>!�d¦)Iu��T�ڜZ.�°�DgS��(t9���J���} \���"��{#_=Sv�$�t�_<"�������ނ��4];8��B�o����+ G�@�?H���i�8��J�}G)��f����,ќP��G@�������xU�ou��D*:�n�SE����I^����m�w^�}��b��5�氈ޥ*�L��W�;r�5�[�G��V�d֕�;=�]'&���l�o���;�{l�a\��t�������Դ}&Q����$9� |��*}��]6�GF��(9�X��nUa��b��Cr��+���4���ɲ+��x���o�\��2�mJg7[E��в�t�j�r	�2R����X��	�@�H*�וNU��q}��ck}�CO�qD�KLD{�>wRN��5e' ��q���r悬�r���W�%ϡշ5�Ɇ5( ��٭�����=Fq���?��<�:?دq"Jh���c�l�v*�%N7W��ݹ���"&|������]�Hp�ϱ�[���[����i<�y�@���g�jɌ�c��k�1,ҕ�t���#i�k�����>�,h�� ����Ļ5ܶ
hO�.�`�yE�O�x)$M7�u
CU �1)��0 �;���Z'E��h�DI�]	$�{�N����	)�����%3��)΃�/��3��U ˧]�a��E��j���S��J�\��KpG�.�x��B�7@�IāXlxVHYEB    3b09     f80��8y�T��
�0�� ����T�r�&""f�0Q��7�<7d�K=T_Zu���H�����"�gj; ��]���q&H�D�Z'���;��bm,D\b=����{$V�'�U���O��{�����^ߓ�@j�`�ЧHReDC�Y*1{h<��;��f�4���+N�\(2aM��@W�ߓt�����'��S0�o.�0)�Hbl\�G@T2���d�l; )j&����z���}/�VϺ���BdQ��?wM��8 Cst��.װB���6�vd�cJ�`��v��_�yU��`��������/�$9 �"�ɿ�/Sl>h;�ŉe݇�A6�����/�f߆$���Za�p����N�ӕ��4m7�hƦ}��X��(v`���凄�Z%ٹ�NG�W��V`&�萜�"P�J_�[<s��iDaD��mk;� ����/��e�CƋ*'�����R���
��3�y?��W4�,>�7�/�$򅎍 Ћ.��7L{T?\�T����D+�f��#rPͷ�N��5������J@�ژ3H�����ʘ���lu�TDi��5X� =9�YN�y�`�6X5艐ޙ}���)OU��Lc�����>���mېj@�+*ir�3�a�&[7�ǎR`���Ȼ�+�`|�����\47��ڌ\ҭYM�E�� �g�����=r��7�G��=]"R,l�&��D ����g�0i+������LsI��Yf\f�)@3��h�څ,v��9#{�x�e:�ޠ�=�$�v{#�|��{g�!E}�*X����
�1Ϧ���3B��I��a���\q�0Y|vO%�������ЀE����G����;�/_B2M�W�H�:yӢ	60��f!�'���<8�ú��*6����)�:�W7m���_��v��.89��E�rXF6�I��t�3���v]��>9�%
x��uѳ#�pqk��;6,hb����)���_y�m7�3ݮ;���Ғ�맸)(����[�s@ʴ�	�>�X�ܤ��R7��\�^%���΁⋸�N����POd�����,EO����R�)��P��pgA���s7�TD��T�F׸�s��z}��X3T�oy��4�b�O�$�
{��eVA���ܒ��82�����e^��L��1J��Uk*���lAn�3��c��5�#А�}\w��Cx�E0%����^�t������<��^G��z�7BV�9P�D_Q;�2�}iD�����A����"¥Bڨt+\�����Y��y�s��3���!5B#���?����y���6��WUfͯ��t�a\�n����?��*��3����X3ם	�rP��,a�W̥�sxp)�J�&��y
���4D26�O�-��A����\��}Ŗ`�"rrЯ��^I�5\(w����-�+���!��s���rW/3�����$�۲`�ƧYJ���M�UqxKD`(nD���w�{���vJ�>nV�����.l\Ag��0r�(�.���h���Z������'�x֑�E�ko�C��+(��t�í	4���[q]��ζZH����V��_�
���3��0�@\Z����H�
�~�<�1����*�&EDab�����]l4s�Tu>i *��̮���-s��d���{c�s49��S�$��zJ�2t$:u�-Z���y�iU��v'm��o�Q�'e�zm��߉��u(v�FTac���Õܙe�����9 ���M�OR/�YF���͒�ރ�<��k�=D葾 y��ղ�+-�0��e��_ �z�v}޹��>���P5�Q[Y=�.�B�t����Z���"�����]�9���j�$�r�?B�������VBZT�k@W���;[І�E���Ԯ�huȉ�p̉;Z��"���^�W�~��Kf��-�AߣHA>�1���fA�3���BY�]����Y�r1P؉��H�^)r<⳴��d� ��f����W�����C������I� |t�6!�Zd�F�/�\%8���:s�Ϻ��j�sS{Л��c�����/F.���G9r��Z�-���e�O���d"_�ss��.��u��DE��8&L	��R���Ae�m-��5<:��3eyBe�&�7<cp=
����P�YXj�K����T;��o9Ws9�d���r����Y�^��J⮆*x�]���U��>�a;L[��'�2�W�R�2)�+m��5�^y�B�<6d�����U���c��@��cY�5�eх�~�Mc^���P�!�[�3߳s)����iQ�1�1X�=�5�N��h�Yz\�����~nǨ��!3UA鮫=q�a# �7��s{C~���;��nOM5��9`3|�E�l�
lY�4o�ZI+�2�H��>�>���n�Ë\#ܓ��z݀3�o�P<a_>��'��B)Wt�XY\M���:���Lŏ�Ŵ�pr���i�A0���^J�J�侹4��������+�����Cl+��F�N�E�UFY��4w$kg���w'�v6#�����^�RLy��� �B������*ڙPMK�8D��*�ozS�`��)�F�_�k�>\���:�-|P�%$ǜ����ɢ���;#�YɭȖ���RH�Á��E��.��R�,٪�޼�o��ey���<��^x�1�������m		��Ky5��8\��ݩ,��A:n'!̾�����C�Id��A����G]��v)-! g�9/�O�i����
xӚw	��"��������y�����2��x`��?�]�r�'��?����LC\y"�����k��VU�4���_���a�%ZV��`x�2I�%�Ɂ���E�LѶR�q��0=�ɧ������`�[�����e j,�#T���H��J˧֡�_�W=�pYK���ʻM�Ba�[�^y�5����5�'�� Nmfř g���%�4�H�+��3J�amc�$5�h���2X�6=�GF sJ�ƉI�H?k��$&ܲ��m�D{�d���|����`^4iMn!�7�/'ZW�Zg!�}b �*غ�&j~�,萒�!�YR�Wi��q'�-��}�����<K�H<H�me�Iv�T��.!�Yh�V��99�d���"k8�5,YT�5"h5�k�.�T�]�G�t_yLz��IZUː���,{G,]a�r�!�#w����F����XA���VV?������E�D�Ǣ�������"(�y���/���x?u���'�}�6t�1`I'<H.��H�\Z��M������X�*#b!����w�ذT�]F=vO̓����o���z%^��`�<>vO��5~#�.+A��s�i�۳a=�E.<���cH�Ħ�Ɣ"n���P�}ˬ�^~�1ư��	��a��p݈��X���ZǦ��l�s�)5�B�M��[��S4�y$�7�kI�B�D�{�D%<���� ��2{���ko���[�T�S�0V+&�dy����R&ND�]���"7V��]4#����ʪ��#�ڸ͠d`(���-�Җ���E����7NA�4�^�x`"�+^�H�y�U_Y����jZk&����5)��+��%�}R&�����PS�ԁ��9I0��%#����[L��u�WUrqu1����"s�>�%{3qQ�ђ�,�b>�'�ky��2��o����RY���n�>�y��Cy+�N;��e��͋���K۷�����kq��{=H��j\\��PJ7W���h������ a�󓱦��0�T��a��:0�y�R�����8�r�u��t �}Siid�E�WBƋ͠�����,H-�m�*O�w'��,���qH�-�va�t�ʝG҂3Fz�ů��`�T�Z�����sXs*�ggq��)�o@