XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���#Z�Tr�z)-���t0��oO<6�����x)�9�x߳0�qN:U��p�,�g捈�۾��!D�5Ź�OBA�H�Za��cbҿH���_�J��S�ʹ�����҇�Y�넜|lq
fO4����F�#9,��㩇 ��Z�c��m&��7�s������ӯ��"��+��˳d�M�{-��v}�+i�e��W���
͊J/p��1	��@'��=�ZF�2���/��Y*�������t/H$2��������֩#H�"�Rܗ���]��#:ʣ��Fx��4ίt�`LZnd��#�ٗ�SxF`��t�y�f����1|ڑ����c�^��g:��e�qxi�/.&��5_�^�˽*ݎc����]�,�`�g��yğ�y�ਸz�UjX�=�527�j3_ņ��yovB�Aj�^G�����|۫��P�D@�q&���5��b\^�o��X�Q�x�+��dEe�	��=���E�>Z��b��ۿ����걔γl)7|� x�C��r'�Þf�Ix�vI�ˁr�j��Y�N�\FȚ��b�*:3�4��H���6��a�r�o�}��|;��d; ��ݗ�U���+X��k躶��$�Wo�mO�(%T5�i�Ȏ�j��%Er?�n�!Ԕ{����VB6�7
�_�Ԡ���QS�	�-.2��w��K�?���~e��E`Fڗ�1YN�صW�g�='8��^���Ǉ<�:��B!��Hv�-���}��XlxVHYEB    5d29    1390
��T��60�.ʭ�q�f�Knr�1 H��Ϥ/`��}�3m-�O/ o��dDݗ1�n#o���l�9:U�L�{��9�x)<�n�6Ǉ�?��T2`��ҀEC϶��#�>�[O$�K�B�����j�x)�k�us�7�o��a�%m�9dL'������U�Ny᲏�N*��&(� :/_/�%��b�*9;�,��b�����ю3��|]IW��� ކX���u�������D�k̋#-�/�T�I���U�5�"3$��;�ԈG}�$�ܼL.e���ĺJ�gTF���빌E�4o�엚�׽۞��7�f���5�Vɿg�00i�6.u�Ȩ|]��6H���T�W,Fr$�p#�Wp�xH`/+
��<�5�S6L��6&	�������=�	�)���[p�$F��^��!��n����Dl�̽��H�9�+r���X7np�r��,H�-!�h;���۾��R�#�d4�T�R�B($�ѻ�B]xlJaV��3��@̋��G�����R|t��70 x�JY"�%A���L�W�՟��\.�x�/8i\݂�i-ڸf>iDF�t��fZA	y�2?�F��q�~��VF�\���n���(���e[��Lg�u�9vԃ�B����b��� &��B���T����845DȑFj�C���Y�kl߳{�Xȉ��6�v&�HZR��%,��N�R����9G���/���R�12MFrC�_E�.7OPdÑQ,ȸ���|� !\_Ug⦾hc�'������GUp��%�I4Y�	�Cz�[fŭ���a�pפ�A���-�*t�iZ�@l{�V@�qf��hQ��oxr���7??�4鰺���7p�2�)�L3��7]"K�7�H�ْӢ0j��]QH�.d�#՞a~M��}��Q��4��u����5�#"�O9���#܊�%�d�3t)MMxb���/�rD,*L��q�t�r��C���q�O�����)�K1ln�߀���/�u2�H]�EK3����@%h]���LБ�7짿mIg��"BN�����
+�&�%҉y�>��W��I�\�v&��!Y�2�O(����F��C�0޸*����*#G�P�*>ם:�@@9Z�����X2.]�.5�����ibc+�ݦ�Mb�"��R	&��fD��T��{��(�#c�1�N���V�����42�)����W��+]��JF��r��������f�D*P�+�k�Vbu�b�+���
ň�<���Q]�-����p�p������ı!����i�Ϊ;ŵ��W�-���R/�A��,H8lhB�~�x8ѣ�^N3�9�?�dS����<�7�#I�\zl��o����X�pWWq�����৷�������5=	N;���$�RD�)�b�ݨ~L���SH7�����-y��.q?�ٞ�f!���D���[�" �WvL����j?�ӤA9�j����U�3{�3�󽽝���c~��Z#�5;~M�f��yx_6��=�/�8��&�l;/0��v�44G����[3�l���K��u��@o|4j~�ᶉCZ�ذ�奰p��7�X��bz�	==C �#Wk\8�òZ�W�	x+������"�B���n�ִ,X���O��nq8�+�O�{ǡ.�`�?�8R��e����Ep�I��5��*��zJp��b�r��2�(��v2��͚W�0
	��i�������&,�{{v ������|�� ���p
8�a�����.�C"�l���\�D��޻jDN�.��tdf;�m�v���c6ʖj32)á�g��*䚴�9/�O�C�^q�i 6���p�Ʌ��5�BA0�����A�� �G���ygޭwe��Z�>RA���3�Lhg<<�#�:�l������c��kf�h�?�D�#J���
Q�˶���e5�	��0n�HI
� ^�pq��7F��X�fHazm�{��f�n�غv���V��-��_j�=����m��^�#�?�	�=*�3�����j{�qJ�04����K�!�(����m�:�mch�
ŌV͸�2�����[dR�D��S�u�u֢�	�t��e	��:�!��6d��}�Q�ѱ�N�F�����ƚ���r��B��1���f�Ƶ�b�o�+	\ȁ���A'H���X���C���ݽ����lƥ.L���>�܄Ȫݿߌ˱~�WW�iCY�B_��iQ�;H˅$�GJ=P�Ұ��ɏ�.1s(��3����<չ�V�<|tQtS��yꂡ����Q�RL#������R�qT�!V�eR�`�Mn��n,L9oQ��mקTB��C�����M�d�C��є�z�|B�}!NN�l,t�s���"T9�h�ʬI?�,�������Z'�E �3���\Ʉ����)��ϟ�GЄ����d	�!'�~��reM��Ԭe,E��U��[/��1TP�[E;޹��r̳K�#���df����Ϋv)v)6{�+8{�˪�f��ea��z��d4�R�γ6Jr���*����k���/����K4��~7zGE)c���8�+kEd���kQO[�ů_�aܹ�^)b"��ը�$D�5�#�i'"����4[�5_���e���0�Y�#h+�W�+sݨ�h������� ���H���Pd�E����EN��8}��T'�+��L������ӡ��wQ�C�'P���Թ�������5���m#@����+��&Z�}ɠ�3����������؀�ǎա�J���h�B
�t�؟o*�s���s�N��Iw-�+;T��f�W=�Z̡5k�w��XC�����`����K�9�d�b�ΣЮ �3%�L�_Ҭi�� ^^w�m��͈���8�������Hی��-�� �S�|�x�>!��i�8 �?�$q��\���i���L�1���3��I^g��A�.0	k�m��ȹ�/Lx@I_(5��*��?v(��Vu����Kҗ͖{��A�*��lJo� )Z�:�vXڦ���ĂY���� �6U- :����%��r�C����!?s��֏��.���}^o�����~���_*����Z�m�`uHV��j{+W֌ d�*@��%2.?Ƞ���7y��W1�o7 ���]����.OC%�F���~�J��g��F�{�d�^��1�4��F��e�����K����ӵo�<��4����7?��ju#
i�G�A[���qhх3�]�:�p�l�ϱ�)������s=�j���'ܧ.�U� Sa#�	a�c\o�=�����������b�y�˔��)1h!�3�s�^Cl��e&��:�@�7�Q�����:��~[3%�t0H"�U��0Qu�r�΅��7�з::=�xԶZ�Rk]��*�+r�[�Δh Xܾ�܍2��"�]z�4��Z��bWni�e&alk�'�-����}-GmD�O�3���� ��r_�[��v���N{(����v�$�u�QF�G���g(�Cˤ��
�0�L���������z8`���S���]@9?<���_����@���6�s�7�����;GDv��_qX�&���6k�a�P@)��zu��R`Ј�7�0��}9?����xbow�uܧ��\t���f�JrV����y}�`0����*b��̈OJtR�(K{Ӡ�t��4j�X�gл�mx�'��A���s`��n��#H��S�T%�����\j�inI��Hv�F#a�
;'S��+�	K	Ամ��*��֞�J���v��C�99Xa��R@�i3��	��qDՅ��A�vf�?�S/Z��4���g��nh�K,�k�u'�]�k0�_90rp�+U��;�>��D���ס�������]Y������~�}�n�\/P6ϭ�^�up?��V�{|�e�����|��z��L�'�g�R��+zSO�,��!'jd\pTV]r�yh�\h^	r�������e�a�ra8��R"�[DE���%�V>�@/�i�>E`)��YՂ/H���Д6�|50�iO�jh��Q�����9,�A}첚xW_���AA����&B�����,*�%Fr跃��C��)-�g�;	�Rq�j�=�� e��-O0���gN�%��@�~�tZ�R��U����Kz�S����	�E��7����&��F���vV�-��	wF;l��X"�H1|A��+��-O�-�|Μ�[�>��{G" hF�Ӣ|+�R��kq�
)F�C!�����61Զ��7D����:�ha��{�b8r�Ϯ/pX��K��7|Q�����s�e�v���������	#!�b��LD{V�mTA�lU�Sr|����)k�+�:⎀�hq�w;H��m���Ԯ���kZV��+"ff��1fض`��̾�����c�x�Q���6�ÓL:��v<O�Wt%7S�9<hǽG�ӯ�;�J�p�҆�@���3n�.ȍ���;A����ʿP��ZI��kI��C��� �xy&� ������
���n��1R~���,����=��SA:H��մ�(`�eH#T�-��NE5����7[�85`C��<���Ro��}c����G�n'ѐ��~k��'�d��K�n�������\a;I�Ư9<r	<@i���GU}nb{(:��G�A`�?�����0	:.��4��xg��.^����}��EMX=��V>Sg�+��6Gx؞L��q��ԡ5�㗺UOF�U7�ֱ©��H�=G���<�%A��z�:r�[2OT.��U�0��,�2L���Už��� �͋U���o����{={�d�GX���-B�]��b
J7@,i�5@Q	ظ�o��a�>-E !Gǫ2�R�δ��6��e�U��(.�N����^���{.��70ұ���ӫ�E��f���X��K��5Ǵ�����)��^�-�b