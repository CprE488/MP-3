XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i��hn�N�^h���G�{彅M���]�l��ٚ)2��:��(q���l�t��[[n��Q[���2�H�ʲY5���c�y�«��+*N�']����Q� z
�L���� I:��p��-�1��?A3��n�u0���}���*�<�cN��8��bP��m0ЁN�V��uZ;c�羁��7�w���� ��B�Z2�D�A�����5l
6��/�2�l}� -�����)%8���Zʹ��.EJn-�g���I�����3iCpԵ-��	&k�y��[J$��fҴ�!국Vz*�	l.8����'bF_
�k�A�V���m񨰑l��',��4N���ٸ���4��K:�*El��ཇ�fN���>�'݈�D�ƀ5�F�9�Ȋ ?N��!@����[�RS�05˲`��}�q��Wo�϶����`%��(��L�*���j�Q�,��\��
�,�2�Q&��-u�f����^�W閤Y���5����4C0&����<�!�^�-T����E�9�B�P��eR�#�ݏ{.l[�`�4�
��d�(e�2s<���[�Pȿy���J43�NT7C��/�m���Vp���7 �:�So���p�C]vS͍�IO�zD\$�KҢ!�?���y$�\�	�����L-~t���On-cY`�ʧ/+�J;�Ͱw�q��s�����ˑ..�FI���!M�+����ǣ;BЖ	f7RO��赡�oh �g��B�8��%W�a$ FTgNܐ�tN���AXlxVHYEB    3fdc    1160�"w�5`����bY�)QҔ~q��J�PН7�r�s}���uӏ�ő�8c,�C��
)�ߵ(|�x�E��n<e.;�KP�OOjP��T件8kk��Z�~\�a03�*�g#l�\���B]*h�'		�>�w��2m�
ȿ("ɰ��L{@��ʎ�)��3����CL��������IK����y��EǄ"��0��{�e˶V�5��IR��(=���h�1Wy�d ���|@tk�=Ե�s�34E�_�:k��(�W��	���g�9|�(7�8�0����%�B�%̿H(��w5s:�2�s��3g�)��9��0�7'5�ɑ۪w���]N����өj6����	i�x�G���l"�K:Ic�T�"7�R���$!jqpk�1✢�0Ȥ�.���ʵ�ٚ��(J�P��.�i�����m��x��)3�<������H��%��f΍�$NFDr���_JCn�Bi�}�|��SS�1d��Az��w+N��_y|���X\�� ��.c�f�gE���J�dE��2THl�#Z�te��<���K�2C�`�
I�[$���0+�|d�-��H���~M ̀W9<���2��
:ڴ�D
~��E)��\��!����߰���CP.N������p�Ur�NߛT{�����F�\�U~��7'�d7DY�N=�E	Q~�������6�7�O���^��A*��0p)_��qN;��IS{�������g)LI%��b�.x^\NH�z�^�a�l!��_x.RՏ�;7���}MXZ��-�fj��o~p8��s��n�z+��ד�
��Y+�9�MP�E���(֡�8�7��V;��`�e��|b��ѹ����˳�E��%v�w��8����Vs����9i�<(���LVt������ ֻ+���{�?X�9�ÅTQ�� M��؃�s�:.�zw,��1��l�~�t��B_v\��Q;\W�H��]��ݿ�|D�)���S�dJ��Jp�(KOa�UO��}�%y6QsB���,}�<��)�Sl���%��*�<��-~�W>tI�_������^�q�^=�rS�(����[���
:j�M��	�,��l5��*H�p�����,�P
�Wͮ�a�
n.�x�M�*��UWn&�A����<;���f	����x�tw��e3D�#зYn_!�;_��	�;9��kNű#:�h� S��֞/�8K��!q��N�@)�<?�����l��K0�����&��� m�r$�G��~�lya�?c����vr+��A�d��HV�ȏnZm!�r�X�̤B�#̈́G[W�s�/�"o�u�B�M���h�Rڒm�v57�7���w���������)c(CT;�w�ީ��x5P+�7B���w���_���},�cēw6&�_�+�v��,/	j�f&S�D��S��D1�h��jyמ;��ĨM�pC	>�ݽYB�3��Il+j��]�5f�<^ST�S(��[��͊o��/�,h���@z�o����#+��DJ^�va ���8:�� hS�\��QE^���=�28��<�M�]��j�z�o�F��&n��LF�S��h�����T�F�N�^����e�c���|�R�ay�z��ͯ�Ǵ�u���;k��;��成������#�Z���G�x,7d*G%��B�Z֓`!��!�S����c�6%J�-�������m�L�� Z�H�e�]�	AZ�ߎH	ɏP\WMH�mJ������b�"��#b�ןiz��_y�x���C�'=��� l�eT�c7`�>��?�§�I����ݝ:n}��b1e(Њ��3�h�S(ռ@��3o���V���K8�&!��E<��i���9��b}h!x<��^�dS;�b��[dZ�`�Ե6�u"�V��P��a5Q�Xk;���3�y+���7Ė�OٺYrA�M��㧒���4mR�+�h����J
� ���|��<��JC	���"{K��������<��΅���$eL�X��p754i�� ��(�8��ԫ�j�Uj -ü�o���R'�ƨ�$D�=�|)mi�A�>I��V�$ܺ�v{o�/�YHs���/����h*�pe��%}�U}�$���J�Fh�68�C��������z9i���5)'��V�����\�^ц����)B3'��x����|�����ԁ��	ړ ;��.?�#4�́]W#�%!�\e�f�G�xf�\�U�s~#F��.,L;*5V�G���+�t�""F���v+[��Al3=u>	t�(��(����k�B$ޓ~d�m��N��%'�c�
�)A�9@�c�=I?���z��B��-�� ���i���O[�,V��՟�ϞR�}�W�����w^A����
�q��z��C y���o����U�r�tD�TmXZv��j���0�q�]��3�tE�>�|�z����W�يǗJjϪ]�H)).�?����6oJ��[0�_>
��������8*X���v��hØ�d�/�N�F��*��Յ�D�Fh�98 J�hHו�D^�ny�6�U������������l%�(J��(	B�h�9��>��ᒄL`�`�@P��Dꛭ-���?��A���$�IT��l#���@�UY$�~��@��Ow���vtu�<L5�����|f��!�Gj-��:z�BeW�z�`����S9�!���:�V[b*��s�Mqw��6^���Wj��$�xf\��2�\V�c���d�����8�:��&C�)z$��v�"���R���2�o��5�c��+=z��5�!� ���X��Fx�SF�?*� OZ�^~]]�]a�(�Z��*Q"ݖ�7a%��ڠQo�>:oCpuxm��}B�Y�4bU�]X��j�����A��=�/�X9_3��!�9��V))�ek$%��&b%�:��s�t�����0cJ���񇦼��� ��uu�#�LʏRt��$s?���:�p.���
Pk���F
�4�K6m���0O3�S�'N�:v����[��K���ϵR�Bqx��3*V=G���l��&1�{��R����$��ׄ����ƙ��T��|�C@�1@�Kf��3+�;���.�7]�Ei\n��UƮr	��[�~e�69|�7�S�w�T��HuUf���O
c�x��-�I�D����z�[@,u��~�T���;}��pPɕ�̡��Q�̵�y�d�|����cɤw�=.���pڅ
A��T��#@�u�x�S�Q��E�o��򛅣��5�ƃ�ĵ9�h%��T�U�).V��D,.*��G5��j��y nb�U�t)�c^���¦k	�8���5X��|�`��W\_�)󆊚;�K�� �H�m:�+[���g�C)����{qަs<C�B���Uj���b�r����8-��&�p�"9�F�?���a�庠|�K*���(�[=>��$���\A�lؾ����'sy�;w��'nkx�a-W~�i9�#c�������3!PrHvc�Fz}�y<�GO�Z�긞3+�m��Wh��BN��w<�v�b���л�˶Yd�N>^v<:�+�j���ӃwJ�|��>��6FO�"��,E�l|c�
c7hm�5+������Ls�[�	�)FT#Ǎ���)$��x�n�6:Ux��8(x��ǓV�=vsj�;
�~��#��u#yx��R�	�9��
u�O�MU>xI#=�S�	�ׯ3�z=�@�z�k>�eQ\�7����x���j�?q%G�&O�'$a�����v��&o-I�]�uNt�\�Abfj��WD�H (Cj�>��q~vaJFe��'vO���dI��T'7�J�wG,�29���tV&	��H�d.Y!I��&����qڙ��7��gEg��W�9+R}x��ݶW %B���K �����Rg�C"g�n�Mt���cR
PX��O���g�NQti@�νÓ�Ѯ4�+�{(Wٸ��\��Y�ce�^���K���M��N��֐;�^���øg�,�\�*R�M��zM����}�5Gh�]=�Z�����;�*uqN������)pU7��^=��u�#v�ϻ!�H�X��mٻu6���t�� ��iہ�d�d|*�?ӧ�儃��,/���&d�<M��v����4�C֪�44N�H�ʉ�Ϊك#do(�p���bn���ΙӞ���)���8�@�S�&�L���"�b-�h��I�'o�`k�	�%Y���/�=]G@Z�����J��S8���A=E;��HbxX.Rh����w�\�b�Z`�^T��C�]�ӹ*�Հ���qGC����9���T�+�����^n�s��mR��D