XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>馘��YH"ұ��m��\����!�G��;w��j�+7���a�
��m�7:�R���dщ|VQ��Tĺ�N�LkU�J@\�B�A�lŽZ�Z�T}�yp ^cL�5���e8d��R��SN立tͣyu&r��#�<�x�����[8M؄yșE��S�{M�fB6�ɣz O��x-&�~�Ҡ�P��B���=T�~�X��D��r�Xz�I�:qo���{ek%��>�S���ʺ�U�q�A���@��y�-D�f�	�p��F�L>�	�/8��pU^o�p�{��	x o�
X5�l��Ϟ�~�h�v�?A{� �~��<�0�b �~�{�*�7�3#�ȅ28����=q�dZ��6���O,�95t\��$��r����#}Ǖ������\�m��u�5X�f�b8�(�6�H5w��D�u��i�y�,���t,�Lg�t�P�WȬ޶��J �Ӻ����P:j��TZ�����&��J�2�/h���d9��,�6��xKA�o]K�@7?x6As�@�f�6�gC��L��␗�Ǳ�p�5�K�~�>�ǉRUQ��7$z-��>������D�$�o��J��rO��Γ�_kT�~{��8���$�ɅĸjMo�wl��'�K��t�ҚY��������0��4�*�e���kc��
��ٍ���V�&�+۞���u#ކLJ�NZ簞@��p]��
y2�E��KZ�r�01W���2RY�I,"�l�w�6W��O��D�-U���p�����:-��XlxVHYEB    1ea4     920Q�@�J���,����3n8�~�i1�����7mg.{��ЩPT�6���=��P��]��j�l��\A��=]�9̉��b�9�fY�m.�j�2��U���̞Ş�� �^G{��Ҵ^xÛ��7w}��QH�W(�N��`iސ�uU��gQ�8����ѷ�x�M�cc~)f"�rw���g�gr�+�?����8�ߤ*�^��Ӓ�|S1L���A����K��A�JY�ǹK�=�9OW��^�59�h�$�0�	s���Ϧ&(���a�W��xb���R�0�%�V02����<a����gQ�Iɮ�*��-�5`�8 �I�V2I�)�lk�!ME�kc�m�W�W�����]��?�4�6R�E4���ty��1}��^����E�9u�-Q�<��&�Ňu�Č�xV���[�>�@
�gv؋�Q`}�m��f����,@(�th��yE��t�/�1?���}j��ʯ�߮!���ҬB�������S+��4�Bp۩HC����]�~�W{jn���.0y�:ۏ� oX3�^2��I���6հӛ)�`�Z��DNq]I���%��^)X`#�&�G!�huz!����k*���B��R׵�w�j��ks~v�����L�|�=^��G�T��e�æ,2
�vc�5���Z�d�l�^d��D.hG�|9K��;s��`�s\��}q���7��5,�������y��\P�Ώ��#�`j2��P�I}����@�ʓ��]���?���* ��֝iX�w�cybyt�\�p�37/y����5�B���dJõ���K�[]�zg^���s��}�f��IW�Q��/�dȶO���V=�!��>�����(��~��i��MF��3���uG!�QjKf�V�$P@�md*��P,KK�k�.�E�OSB��q7
�Ri�.녱�_=��+��ʑ�l��Ym��
���MP�|��ؽ:�s�\�hu�Ũ��b	�6����(����֮'=���0o�>V�*�O�Z�O��e�u.��4��I�3���F��+��c�	[�����
�PB=�� &�n�W[��ĤZ�ȑ׃"I�c����S��.)�/utqT��vڮ���yG�N࣊�B��G��(���qq�p)�ƗvĻA�b��v����nFi��D6�S���oo�_�P��U�,y�4 ��?���%�Li�ڮo�Ԁ鎲�>�n*˺Y�$�ys��3�@
Q����6%�TQ���Q?���?"�۸v��<��`�G>L��$U���#� =!�1j�b�x����-(#P�C�J �<��vUK�%w����]��q!CҊ�>*:�&O��ByO���Sg&$��
V���fUt�z����z��T�+�#��Ҏ3	�Q��<�:v���<rx�ָr�3Ω3s���!�.q�|	G�8�B��r�)uȥxZH�ٙ*O�e2D�d��A���O���s�d�?OV	0r8l���S.�������q��ݺ��CZ<�::������c�D�Ƕ)�"�yݲ�?DsL�@bpH�F޿��#]y��-Ϯ���i��U��k#�-�n�0�$���a%v=�p;� ْ�mK�E�x^|�Y�1����{���>Y_�����#R�m)�z�{��νj���ʾCon�H�[ |�.(���>>^-2I�
`�%	�
4�@:��M��~�����n��%'[�-��JL��TG�0,6��D�U��x2=��.'�Tr{`���WږB*�1�d0��{x����:��M*��w����D�a�K��'��L��yl��Ov�������G�x��/�[�p��-EJN�>��� � �E m�u0�F��+������
�E��qH�J0�0��+���M��&��J7��4JT�S+�o	��,���H���Á�����R�^'�� 4��چ���Wa˗Pw�U.�#!*��m�HpБ`;# �K�1Y.D�.�����;�F5���>������p�D$�[�����=�A�@�_�D��I!�*0/�I���4�*��<��sGL2�V�3vJ(YX���{~���Ѯ�3(���!$=�*�w/�q��,W[�Nfxw��4�M��@�U��r͠�A��y��VۡT��*ٴ\᧪t�Ob��,kKF�`-H�4������a�3����MN<9�H�럂H2�`1�j!;҅�券;���zp���Z��k���f��e�)H~0�=� Hh��Tx�G7$^�-Zؚ��d3��A�[tW�_�25G`*�Sa����>?p�˿H3�{ �*�r���眊��