XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z�惚�e=@���A1�X�Rȹ�|~e-�Ԩ�''�;� ��)�6�YZ5#�Z3̘íi]]����1�p�%�$*�iZr�<�[,�'��	�qg�%�AHm��[�pSPnyL���*ܱ* @���*
�D�"/���l����K��8���y5���8����htM�$��������,��M��;��j~猓��d�tz���5+l�m��R�WY����`��7��l�j�5�d�;��ܯ��9ʖ�4\���"�E�K�~+���� ���n��#�NȮ���m�Z��D ��
�����)�@��0�xC�������wx��u��{�W���?S'5�yH�pA�T���F#�����v��F�x��}V(���"�+J�\V,a�30��:�} BA�M�C�D? ��ʥ��TɈކ���ϣ��4�N�$q��G����ݐ5��VzҐ�<��-Cg�� ~R�SzN&H�ӓ
��_s;��+�l�&���a�yEV��8D��I�p�h����ʁ��X���o��6��[a]^��%��U�K��.���y@��q� �ߊs��'�������������U{���^������ZaJ��~�u;WK�-m�_�]��ڬ�H7��.��`���)���j���Q�*��Z�R����$� P9�Z�h��g>�]8'NsR8�6�XX��b��S�7f�t�Y7��ڐU	D��rJ��5�����]�>�\����1� XlxVHYEB    17b2     880DE1��W��m̈�VR�D��R�S��}E9�	���դ�0 ��P�O��(�`�����~�+�S�V��	@qJ;�=�/b�t��4���*�Y�3�_��+�(�͈/ʨm��'~]7U��u���e@�u��)��;O��ª�0��D�M��w��:�0�5�-��������K��b���ϞȴT�&G/?9mӏ��x�k��vsIy,�$f9<6=-���xS~̻ʝK�r�!���&H��'�4aW�s��ER�k�`��W�cߨ�c��R����5w�TAj__�M5�:UT�����|(l:!r,6�'e3��r$�s�$vsAP:'��`��`��̛Z�ߞ+b��;�[�Q���x�Ls�[<Q�H��p�>v2��[6���L�����v��x�n�z�fـ���^��mcν'<5����H"�i�g����C'�EdL�4���k��t��C`�� �O��/�R� h�ݰb���w���[�Z�����-\-�ȯ:3����4��_�^�y�,�2mu��g����牗 �c ��+��숝4�4£�8�$�L�&sp�
�9յ�e�,E��Q_,���J��dy�{�%��q��v�z��|<UY�Y����l��%x`�Z���<'r�E���Y�Km �]�,��ʖA��G�u毕��x�����p3	�>~��i�.kL]��y|H������K�=������� �Z?e�����C������>�|�&O�
�^�+�ʕ�"2Z��<�K�=N{�Y@�鋩���Fyz��g=SG��� �	$n*��cm>h�W, Ǔ�)A�}�E�>��T)DB�F�B�@�4�j��*95����Ez�����(��C{f?����-G��i2E0�U��T�Ga�0[F�	'$u�A��THf ��o�cV�ti���O��k4��*�&s����";�6^T�Q`w)�%����n�LZ�ADH1�~ {�T隮��&���L+��BR� %��7�Q	�q�$@�u�P�c�[P��Z0�ϳ�r1m�K;,m-���Y����N����#��z=u�,�Y}�>H�+���۪N�84�����H��Ռ�򣁒r0�p� ϊ��[w�����&&�p*ş�}���\��#�~zf�_h!�b}�����t��}r�- M�m)Ȟ�*�|7y�/��_����Է8h.Kdc�T�Y�i���B+����iR�x���3��i�z[E��MZ[�\�Brt��`�5��t3JXS�I�0�vҽ��
��[dD���a5�@���;4Y�rIs���ܶ9��pi�>s��W�\���{F!&R�x��8IH��ŏcnغRg��|A�a���O���YTR�������ӧTHD��F�R���1Eh��] ����[ZW��m�'�2�G�z#�	8&S^QUP*��ONP����*ٖ����x��EC�%�a�����~t�R��w*B� �� ���l
��D��h�vՈD�nvZ�\��֤7���h��4��z'�\c�n�zPj~t�I�m=l#��K�E4'���N�P�+_�C��*p�D����h����hc�jpC�9*��|�K����25|�D�CA�P���(QՆ�����6��#� ���iZ��U���<◰�͊����/��c�-�epڄ��!U2�������`�I~�ϙ���ė����]�_���T⊞0�@,1��cZ�5���,2Α@F M��횧��+e���ߚ�ׅ���-J��bT�Ε��i���E�\l�G�t�\�E������j��=�շ�Nf8��j��y"�Na�&CמH��4�X�IC�D`�����1�]�©��\��,z%�{�b6����O�R��L�f�F���{^ZcwNihR̠��/�ȟ��w��#��%ꄜ	˩(/�T��3�����(ϻ��{"7Ƴ�<&�L'�#�U y�|�2@^�H��T���"I����w&�G�R�KJ���Ƀu�*��иjYˇX�@���C!c��X灂7���f0zx�'):�����QH�RK��a�x�0�A�^��z�T�su�jTm�qCݞ�A��C|Ȏ[��h���ܹS�#���ӈW�x^\��6��B8x���N.t�c���G9��