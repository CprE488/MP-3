XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ຂ��t/�I�D�vH����;���@\�G��2��j����X�V�Z2��e�=�S�K��U�M�=s��n����s�E���E�n�ZR��̓r�9�sfHq��eLmT��<�Y%���΍�
�T�����C��8���1��n/=��qgt5'����=��2L}.�*�p��TB��[�ǜ������ �n��N���H���P��PQE�k�\��α�j�i����U@'x���y�е_�U1�{��Ȱ����E��W��8���
��^��҇,$���]�B 3�;�<3 �=�r�<@ 䐖�;6<\�2���1�k��{�TL4�4:��R�Xx+�T_�����_�X�[sB��Cȼ*��*��D��/���G��k$B$ũGA@��,�
gB^B��/�>�#y�E�/���j��d���m��:"�&S��X�&��ax��Ǘ�i�i�b�|��.��7EU��ë���A��*2��#pb5��R�9�w9q��Ok����!А+~��ƳŽ�Ğ@�~�Vp-x��)VM�l�P���L���$��n�UX�"�eVH��a�f�ڰQeIL.q�?+u?5*�� z��d;��G�)ӻн���h�>b�˵F-K����������M�(��� h�ݞ4�N��X�R�i�J�N9p���.�fm>*�K�X'�K�o�������7�����5	���� �	)�Ky8#����)��jT�I�(��0"�V�".YB���.@�RS	�s�E�?��[�GRY�XlxVHYEB    13ba     770K�!���`H����`�L�.#i���"՟����U{���(��PI��V��� j�
�o^�D_N�,h!Bɰٞ`w�f SAIgI�} ��@_'D�������K|"=d�3l�qP�x�x�K�w�`=nN)������@�L��gO�
3 �l�iT��P���g[�Gi?ք ֺ��h �P��R)�SG�P>qJ ������J�8'�Z>���R"5�s����p����+��(�ɉ�T��@�s����3y��1��@4����Yc��R@�p�_�$;�������h.o���	�whɴ��š��\|���^Fv��$�[`k�\��H��
����7A2-4a���v�F��*xu��:�����Xj�O�رc"��Wa����q��jO4���78o
h�?[�?����}���b���Pl�@ >5^�hJ�� L�4Qt���#'�Ɨ���C��a�D�	��H�C3������I�P"ܬ�ԋ��r�s^^8"c��&�(��'�X��4��P����8F�vMMy	�h0;K/
���Eg�D4ZJ ōHQ*�s��A(Y������3����7COI�.����%����xREg�S���CE.�߄W���a(lԠ���"����4E3{��z�e�D[���Hd�]��ɳ$]��,�g�N��뜔�,F�
�߽�f8M<,�9W���,B$�;���5�������<���������qA��;�9Z�0r;���RWͿ�Q�鎏K�m�';ku���J�%[�����r%C�2��)����e�;��Z֐J�eI��pU�/�g>Ss`P�]�LR���[8gr2������8�<�HBR�F���O�5^)6:�팚D�~��p��V-jv����;s�V#}�+�䞤��� o�:��w���#��ݐ �;HE�=���p(g��������~�ɝ.}�ao,��h2gv���_�������j8��fJ��ϧ��O�a{ǅ�!W[�3R�R��Ӕ񱇖-gqZ��Ľ)�$��;�"\�5�c.�W^��[9�C�#�S�F*=�����ve�j����m�����S�qh�"nw�i�i��	�(Ks��#�����Z�[_���ğoB�d�L��M+p�|%G���(���a}lp7��RiaU���I�A�㷟h��d���3B<����P6�׍8^N������ٸ�	@\�k	:ߩ��l�ǝ���vz���^�/xW�}���-�t��/2c�D3��#H#bڔ���ų���du<�@9�u�������t��d�	8�\z�p�Ou{�;����-9���̶�
ȁ{O�h�w��Qf��
���<g�L��j�0�.[\+��
I�<�Ug�!Ӑ�1�gJS���Ug��31�c�R�7��+Rj�{�SQ@�*�A�M �hD'��>l����xhǵotz�?�K��㩞�����s���@K��g�����|!Iz��j�V�ЙV?��}��A">\���2�.� ����[-����n,��Z`����W5Íz�C7����{��8Ӄ$����PO̧+�w�h��'�����#vuպ;���õ,=���fݪE�\	�	I�\-\B�D� .
��q]�׳?��R���ѫh�����+�B���{��9%3n�յ<���bw���U&��%���܁�R�d�ܷ�����!R�:��&1�e��i�KM
�o��o,��+ڻ���? ;.uж��U��%���(:#s�Ԗ���v�/��	���.�ճ�����[��dǦ��7M�� �l�"����E�q��?��AB�WQܴԼ �8��m�Q?y�
\D{[