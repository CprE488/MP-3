XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`o�N��;�AU�?��W{]k}���X�������;$�8�?���ӴS�0�̆����D�^,�E����-���lq��[�	������0:!�Ҿ��m�������J\[,��g�ɉ,�	�.b�G�O�ߦ�,��F&EKǜ���.	�.jo��o��<�� T������������c��\�,���I��|�|K�_m_p�d�\�~e �v�G�)��W�5G���3oסcd/Q�8գ"�4%/�Pj� U��Ճ�a�(�'׈�ш��R
�L����1�A"E�-/8'��W�s�w�:��U����mQ\�;�b�4.	k[@�y�����O\�/�\!�y��d����֖�fԥ��?X_8!v:�RyE�D��.vK�O�[�x^�c�ݯ���A�A� ��:Ì-]M	2�do�4c��WV�?<�Ki��'�j.����Sob{G���ï��Q����2<��Sh�
�Մ	���]ɪ$\�/s��tJ��H͝;�f~EV�ʣ�K�1��Ը�3����y�>Zh=�^�G?=����E3�(��+�|�dT���/!y:&`��
��a	�|����7$u!�B{C�L]W���ׄ#zA��<^����DC�D���m���?Fˉ ��d�ǩ��$s�;�,smd��;��p�2�ht�z�Z%B��g�W!۹�@�}لx Ӧ%·�v��r�����AS�n.M?��(�����1��yd0�랇��FS+��/۟��W/���$����XlxVHYEB    925c    1a60�2oU"�%�q�H�{W,&&�3����	8����t��;�g �����N��LzFΩ�9�U��I�@���7�
�����F����MBa�_�yq|�\
�I��~��S$��O�y�{��GH���q��H���s�ab|�6��K~� B[���Gu �^7��B4jgq��|<;[�#�	p]he���np��Ʌ��Sժ'�jd��1��0l���H��l��4������~��6���~L�o,��2K�+���҂�X�]�,CDeO43W��op<ۗ��h��4��N	�ԃ{Z��7U?��ѓH�#� [��;��m$��ǝa�KO�b�B���㯷(��qݬ��2^,Px�����O��TA��]��<4��ĩr�i��.�K���	�9	���zb}lKu|�Y��1s� �N��8�����´Ȑ�u��ЈuZ?�FV��w"�����aP@�����	h�P�]�^��{`�0~t=H0z�:�ZǹJj�����7��B �������@q�*mp�U������Tu���É�F�U����u`�LY��R<�F�`��H߫�q@�^�F����s#����Lb&]mԎ"{��I�l}�GD�O>���ڷN5ē��z���m'~��%Ep�M���6��dA���h� g}�<�6�;Ơ�!C�aF����h���^�脫%��7����^6J��%^0s=�-3Y���ll�A�tN���U���6N���|�1���Kʝ�@��f+��O>ޖ�,iGP���v��vLDCr����c����dR��h�{+CF�S�q����I:�g��>t�]�tç۶h��(Q���up�}qfn9L���3�~��4�0��l	~�d�M��DG8
�>�u�n��	����pj���a Y�}NR�hN����Z�D�[�٥��r��|��ͤQjs6�|�C�f��b�Z��-&C����1���Ӧl�&�ԕ_�5��Y$
��4"���P7��9��ɽ�ZW���i��z����l��o����XߒM׏#J�9�!=��s�Ew�r�����)�Rwkfw��$^��ȓ���B��n�A���契7�Ųό���[Y˦z_F=p�ɻ��T�Û�K������j��-6�B����?j\�W\|�ZAY��U�]D�6�[����U"`vm��E;a�SPB�Z�dQ������u�i�����o,����"����:�I��f�����Y༙h�m���z����_��A�KɑH�����|V���C]��[ fo�fd�����}��}���"�z�6m�v�v;����%�q0?��i��0�o�\beť�z����d!�e��s<�m�"w0�kt|N	4{�v_BD� �����d�k��N
�d^^)P��<�zћ��6�A���v�a�����!D�(��Lݾ�Ko-t�����psh�}o)?w����,&7����?�p��#/eK�k��j�}�x4W.9��4�ԅ��(L_�1���sZ���
��U,�i�pB�ޘ+�n�lmL&�)&��-�v��^� 9[��7����Z^�p8��W��I^Z]�|2���]±:���3�"���m���"$�@"O3��::��)$�	�0�E����>�a��'���_j8&|Rl)\�[F#s,S]Ӣ�kg2���^RLP8vգX5�zLzI#�	��{�7Y���!5���pl��s�a���}����ǹ�_�j�42N�PG�����K���W�]8y��D�h�*]3h�y�������('��b�/�ŀ�m�K�X�M,��=�%�ѐ�������EYo�@�.ݳ��zf*pRuֆ�$c�cO�����r����ru�/z�C�xh�#�K�
�Qq��+��G�w�|oX3+n��p�?(�G�
�����)ek@���O�2
���� �:�pr��8�?�uDU,z����[6{���R~b������ֲ�ڀFr�I9d��[V��o"��Im؋�Vd���/�Z��}��f>����3ZEt>��\)|<&�S�6K���8?	{56�	s��'�Ut((�F����.�s������s+��/֪3- L�8�MMy�m.�,��+������Q[$t�L�����Ϊ輵I]������}���㚪�E�yY�/����5d����'I`,�,g������?��jZ�^`�t+Mx���(��h�n80������V	1��!f`�h��1��w�Bgr=\��$�F?��F2tzC����r�~��i��Kb��<O�*yI��;��&boE5�= �lOګnm���T���&{��< ���8(��p�SB����.3Z�L���4��9�r��Wp���]_n��Tڧ3��D2kF!@�������З�J�WtMk2�������1Mx���`FȨx�?��rS�'*��$X���du��Ob[�́9�ss6���`��p�k�8E;�.�=*��\^m<nU�|ڝD��5�5�Gy��VV��DA���g=�v�\�yi7m�9,,����s��7�_R^齀^�J+8��=	�xӁDs�B���������"�m/�����3~ $���k�^I5��S(
	���wz��9̉ړ"D�?����L����QhxZ;-��b���xTN���y�*�d�"�{��Bf�����:+���9�;H����N�)�tO˃����G*�Kt�=��
����uKe�.E d;��Eݑ�h�c���:<����VRVN#9��(sϥ�� &ƳF㯚���p�HC��r̫�Ǩ3�@2W�;�8��Fő�k�����&FwhA*��> �7o	���+��g,���L�����ĉ ��+bM��gC�5yM���`�v�;�m����oH��أ�A&�8�m	@�%�BZ
#!��g�j9�$��	z��!у�f��^�=�H>7������K!�Qr%S�k�:P��w�!�_ԝ��w��C�QM���T�#'C�<h�?�0�X���1��D���ꤳ1�R�»�^H �ׁ�L�S,��j�B�>?I����U�0Ms��%�\�*���,�����>��욇�X_�åf���s��g�\�A�E6G`$-�4��Z��a9÷N|�����NA`�#���80�1�!y�oY���霱#c�"�7�|�+H����o ���y������}�x�]�A�"MV��P�O��������.���p&���Ug�����Ѻ��?<T�l�w���GB�j��J�R6�K*Ǎ� 18�����r�5R�9�.m����dm%Hd������Wl����)�������n�7�G"6�Ǡ�Lm������U�^�r�C]VhU�
��ocKz��^�"�Y��S0O�tB���k����̂.��m)U��Ct�Lj���`�i�B>�o��2;v:�,��0����7�JKd����`�y�].E�:ƀ�"\���lPI�T�R���T0#!��� f
�k�~���q���ӘjRH��ߧzAKvcY9'6�1�Q�V�� ���W�������ݒs?{`,#<��AKJ��r}�(�X�>i
g �OM宦���)'�z�
T���p�dM�Xk���'�X9�����/�\�SV&�oT�Ʈ��h� "�M���8���;2W^�����Ǉ��Ytb�IB�4�b�&��l"B�v=�|@�(�2����p���L�s*#{?�����#���MujIB@��<�c��gn�\��}"P�,���<�s6�Mɖ	�v/� �G�Y�	]�i�ĭbP�o��.����ƮY9>r�A8l�z��V��	��q��X��.`�D��n6�vW�X�Ȏ0<���C�!��>�W������m׎	YԎ��&MڎF?�T�>���|�!���K>(HpxP��whD���������N�*Zˇ �~�ԁë���`�_+}W�醊�K$.!�?��0��O{�tK�\�M{$�zO�O0���^��\��XQ�8���[�H~�*���(=z� z���`�7����8��<PL$]�ǻ&�ԝ=K��0ί��a:0��_?�-G\��$/R�n�'�(\�+.qC�J��ھ�*��r8���G�J_�=�"�Z���
?��RV{z��t�7�6�uGU��I.?gmyM|�	��L�Y�{I�{������~�[�ܣ�$�8��H��" �R��%N3wP������9�r�XZ�ȇ
��g��G��rQ�������X;iBpI}�_u(V��j���>:i�>�|w������/�TCg�uvZ�;\��k���}���H��s)���u�c�Z��iq'{3���Z.�a谯H��a���$�B�=G7�����6�(�,�c+���ۦ���R���;�޵�|u���@cOC�~�L��.�]�Zr3'�\mh�T�+��K�����p)���3?3F�TX B���8���&�����
��;�g��`AΆ��������D�.�8'�W:J��]܄�����h���0T`��q���"�a�j�{2�(���B�B�-	����sfm���.�aW��=�F��%��g���%�- )����@Ob�	�JҲye���o�=�Ƃ*��ї�K�d��ňkp�x�c4�/��~4V�nj2�͢���I�|y�u
U�]L��;�)�ؾ����&�3-��%��8&� 	����P��Ǘ��m���p�����q�qr[�+�/�R�Ԕ�,�$ɇ��v���1�>t�Zo٦�M�~�% j��[�����ֹj3T���*p�LfN����kn�Ȝ�=zj�S�d�BJ��vYt"sO��ޤW.Qk�"����,��f,�U+gǙO�^���O%�����:�)���w�=��=Pˁ���v0�ּ��Gqaj0u�WO1��/�=�~�;��g��&���|7J����̧f՛��Z��{@(�%��5�C�Y�"Jc, Gg㩓�f�8=��"8���������@�oI�>r��O/~��ߏR������GyJ7G����6�����7J�׳��^|r@�A�-}JP��t����d��P����-J���j��(y�o�> @�v�o�?^C��ܘ��w��8e
kBW}++�|�>�F���v���6���wo��w�m6.�gWOD��˅"��S݅d��ҿ̀j��
-<晢���ʗ�#��{�Z�3v�v@H!�b����E��}n-��]�(�Prf��絬6-��\����|�D�63�F1�'0���@��ǆ�� B��,�_�`�������B䴮x�c�+LUC������m�w��22�j� Y~`u��M����;��ҜG%��Α<��/����5u[ |��G��xC��n��Ϋ��QplRc�r-ܚ�Wz%���"(�8�G��~����Lt/S��H`�av�_t�4;b�q���`���b)_t��S������/� �`+tTy;ҥ��7'��4�M&^��} @���?N.�z�:�x�o'��Cc&m����獫�,J&��^#'�ҍ稪߫�\��&�NK�-�ާ�@���W�ۅqU��.�T �H��^�m@`�H۱�OշwT�%�3ޔ�����������!�hC'�T������:XE�(��1IZ�~���ϳ���M�ŲO�?A� (�EA�م+��?��
����sļ�+�E��j��� �����go��E�����l����f��Q�Ci� 6��%� �)�H��7��x��RkD��&w��S*���3� �!�4�l�ͮbϢ��E;��G��������8�����DR������1�
DW�d�tCV�\��$IX�c����*�������je�����ޭ|Fנו���6t֌��*�_�7��w����� ���	�J��aeqށ�m���Ak��q�y�MN*J߈�����+nw�j1�����N:�LՂ��:f7���ھ���p{��u�6a}i��!p���},�)�qM���6%��B3����Po��>�v���<�L/C�ۦB�vU�t}�w&ai�CҫT�7�i$����JU�By��k�삯A����N�cJ<�PE�߬�rH��"�D���ٺZ�^W�q���q�b%E\Q��NPдM��~���LCel�˽�"+>kJD���)���/�2  �Ѷ�XS�&�Af�<ґ�Ԕ����'j��Z�B�|kt�P&ގJw��Gp�=&2L�vE\ߵ�N�}Jc%�uk��N���0[e��=�R��+4���(��v��P���52�2wc"�{�%@hPn�' ��nX��m/fs�~�އ�;��(�/bW��q��:	�w�e0Ι�2w�o2Z����.;��O��[��\H�Q�f��_ �{�
<�'F�d���\��P���b��3�$���5���o�x��5�Eʕ�����<y;a�6�	���*�F]�����Ԙ���.��Ey�#mO��B5�TY���m$�m(���A��x��ֶG�-#*K�3�l��&���n�C7���3���r!7�ֲ�[bQƿ���/N<���86T3��>X��Oҥw"]��Y