XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~DD��Y�%�y�2-i��(O�3Cޱ$����m�M^�BIZ��� S:���K��/��k+�=,���oQ0x:�Ϙ�=�U�����X$���e����^�C��M3¤_&�muūz�F~�EеH����l�(Ð@>�3F�wKyQm�����~��h�)�)�{�[Z��%�=�g���+�z��=O�V�x!� ښu%�t�c�g������t/�Q�khL!�B����QTG��N�xޑ��(��#��V;�S@+���S;��3@C�L��|�����͋ԡ�ª�Oc��ʚ�����@� �Xڄ�e��MK�@<�@���4��[��eN����@���"�6�Gr9rK>F�]�H-��h�\��q	���ʀMl-�,}1R�s�tHK.X՜�4[�p���<�^�M��M�}�gYRu,��Jt(���(,�������r;�~F`��[�����Ã��\�m���w��*�|��|c��:�����p��v^,�k;��*y�C_�	�p9�Ix�*�A8~�~�� ֑���6�aU�� 9c܇��s��g�mc��d!r�e?l�I�B1p"��3���X�K<��`����J&{�����ƽ7h��(����q�����,�]�F��cY���ҧ�A˒�H#��h���x~F�{�*�`�Lq:�6�����Ns0(&hE<#�F���}>���	�L�[�w�҉��&�!%�ж�n��\At.n�Ï��z4q�hbR�pXlxVHYEB    3d1e     fa0	>\�oÞ���ǚl���Z�_%xnN^Yمn���� �S"/��N�mʦ�W?6��z9��/sCDk?Pn��kz�G�f��d/q���m[�/١C�8��|�S���'�G~IQ��N���H�~�]��[��c�I�+�����C�>Ӂ���k����?�Y	[�W�����
�O�#�p}��wh�����'�(q?`����9ll%��v��s��Go4q��2�|�
-ru�c��dM<�F�N >�h��(R��a����s�'<�i�d��!D{��)������vl�@5�k�)��pƂ%�T�	੄�`�U���7KK鹿X��ܻk���{�'kպ�m��Rx\�y�����\x����y�q�vpecf���8|/bվ��1�l7�$:����&�qa�ε���f�{�s��a,Z;$=�� |�Z*U�Zyq�A;0mk�3%�'.��k<���5�\P �M�ᡙ��� �FM�n�w��^C�/�������w1=������)/oK6���ޚ5�[�[
]���VoCd5P(\���#ګzA?!�*��������3��aT8�]��H��N�ٿ\�O�M��D���$�R֢����`����T���y5*��7�_/������p�s.����N���U��F�q�Mm�bl�����?j��@9ˢ۔2�"�ǩ���sXf��kF��lP`VB�����E1�`6;P��'8�+�p�r�#��mG�����i\��0Z'h���=.����V�=�;�N���:3��w+��PTN���zgnY����w��b���>���9����`i�������t��j�@�6���%X�lG�,7�t���Ѻ�
�~ŦZ���ޠ��������|AA�2�<Z��i��X�{{�h\�'���rC�������,^�}�ds�G-��̶02��q7�~���2��f<�/
�n�����~
%�z����Q\e�i��_)M=����0V����#΄����{�J[Hc�E9DC��As瞒'oz�����G�c��������� 0ɝ��I�6mݱO�s�)�&��tk�T�j�s՛������:)�Vg.����ɉ�Z��lI�b[��DV��@I׹�摰(`��&U�T��J~�8��9�N�'�P�<��K�(��I��l�4�By����wu18��r� e2�MU(x������7���;��2s{`G&�zu3rX�W�2�N���QJ˟���"��*��__T�)vO��ue:�+��|�ÅQ�>�%�	]���B�-i�1����y�R�7[+A�هm��-n@�ߊĳ��������g�8��M�6�����I�Y�I�o��	'Ҭ�?u���;�Xr�����9&D����o��]�:�f𤳹�N=%�BW������DL+���;��J��m�g���=�RtA��ͼr 0u w/G�Hn	����_�C���D@�w����[��[;]V4I����f�`0�^2�]�u�a�]�J�N9��Y�/����D{p(��k������k���� �r�y�1Ew"� Ii�a����똍x��%�A�$��H'W�yv�y��\8��q.��n�#mo|S���~~iR��3��л��=l�?������ǖJW���0��<�������
������@�v,)d�*�s��ǆ���>N�	E�$��W ,?[���D�`����9�} �ɩ^6w��Z��H���f\��D��6ӜYc�U�#�|b��E�%4	���l�dnx�:��m��F��D��Ry�L��$�<#������mZv��� EqBZeq|qQ/��6�?�=|C��r�P��Dj��%���-��������8L���9�47���A��1��;ۋp��Ç�&���csfވ��]X���_Z��J�oz,�ڕ���pK'ӛ0��?��io` �"S�`l�v�l���:�UG����~]�;R�a�?I.�n����\@����w��t���c�%k�Rg�g=����VC��Q�w��vA���F�qǿs�a�4�N�+o=�&�B��9!F�|�`�v�e1a�G��B �f�����GM���o��X8VW�>Ⱥ�����hA��Q���Z-��hV����>}�6����+#���#d�a��������e�7=�������ve�?���%j`�C�\N4����F�#OO�>V�X ?4O	���� �W�XČ囐��)���(���)��d��x�!��i{幡z�����}���vm�ܠ����o's�+ǘm��@鱴6�BSE���S���u��J�_E�6��H�I�o�j��c��R��"*��(=8���Lb$i�?׵������ΰ�V�G�&!O�+-�d�<��}H�	�'*r�á���|.C���PL�g�����'�/�}��
������V�S}�^���\�C蒝:�F��'�׍B%
�5a[��)��"�=D�Y��$�0�.��'�eQ�xrQy5�v~H�i;�Qb8�;RXW)@|��D;��8َ9�;���	Z\פ�aU@��+TĴ����pR΄e��h�#[�,��v[C�������c/�pe�|<��ᢳ�%󲜌���3)i���F�𥽶�M�1���!���8��S�<l�O�rTV�*�G�b̽�
-!TrX����5��
�|D�2SMGo�9b7�mwg��k8���kdTИ�m�*�E�+Ok>a:6�r���(�(���-"+��- :ncc��aB#�Y��`lX
��+�
���U�����0�~�fuN�A����=j��	yB��}Y/�k�U'�����WY� ([r����C�Yj�E���ދ;m��|�uǠNW������~� �.Z��kc�5a6��h}"�@�ߠA�b���K VG���p��e�Z��^-�=�-�-�v("LZN��0��n�R�����lc�\���Y9��LM4%�XU���{�8�`�� ~�4�w���1]R!��E�z�,��"ў6{
��<�]ɠӵ�V�#M��7�-�rXT�U��a�� ŞL�<��\��Ly.gߵ�l*�`��/�il ����1ހ�L�>�T����Ui��zd���#�3��?�{�th;�ތ����i����+�j���Dey�M��r��;4�1�QO�*z�$��J�ȧ��E]�^��(��.N�b����q���P+5�͏6��B'h�����ڵec%>�t���8�Ԍv�6/}��s �ᓞ���~LC@�|i�n����G<v�ĵ�$!F'$t.��^PV�l�SxX�}�MΜ
zjU�����ud�8���.}�@�&t���;�n��s�����"><|�v<0��Ϗ��?EW�_(����K0�B��u\Ɠ_xFf(��D?���<��
����!o�`\��Ś^�7������>.D�w��΢������������OM�%X�����GPso
>�n�H�Jm>LRY:yW�jQ��I���IL��dY����֒�5�B�Clf����k;0���� �aڔ��A#�eAha�wԃW�f�v��W:�I�UI*#_���
ʲ~�o�<tn��ݓ���^3ü{���GD���־��V��<��4�H�B��^=NvN96&����~� �ټ�$,�=������J��&%��r������`ɝ����E6��HE;6f? ��e��p����Hfp��Lo�T
Pvp3́��6c�#B�"&\ɳvO�.����W�əX(K���U91��D4F����������j�.�b)��{P:W/O:/�2A٪�w8n��ya�߃w��g*�Ox?]b���0q���F��s��P�̾roWj]�ƴ�~@�%Eԯ