XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��CL�^��;��F��t1PV|i	c�/h9\��`�5���r�Lk�����������o�������ࡄ_t�����BL�kbt�Ow�3���;��*(�Yl؍��gR���]��j|<�9��������@R���I
^]�:YJiGCC��upa�ߤ�Y��Us��7��0�k���g�#�rP#y趇N��!�]������G� nu|�o��o�7�ZG�C�z��3�~�W����؍3�ǆc�����B��EN>���K��g�����~�;a��H���~�����޸?�3��?\;]l�K�3m���]�.� �|@7����|�6���B��Ap@��J�s���X9�ˁQ���<���p7�vzA]�r�Y���Ć��V�W�nO�鋩�Q��{C�g�Dօ��a��)�:K���%{�ؿsQ��p����Ǘ�C'���T[;}�X�;,G�"�avj(�����&��V1�m촑Ƶ$=C���ShwD^�%;����=�*��F6?q�e:6ۋ�*�=l��(��r	���/�]�=崅��J�c�1*J���1����^?����SLf�h�L�_u}���Jp)��VǇ���@��L�<�2� �������v�i�z�lM01��l��ILo�E�6΢��+x��� el���"Ë�/:}�}N��`Z�����m1D�ɣ�(q��x����V��G��:��#�����'V�as�*�.<#e�U Lk�\�#�L�([�n⌁^��XlxVHYEB    70a6     b90�B}��[��r��)��7�M�擴��/=w�ը�V�]�\X��f9�ܳ�)kI/\�$��wK���U��NBj�n�C-y �KAu~�AL�{Zǣ%F[	���X�s2}�4�҈��1�H}�W��T,PR���a�+�\��.�@�F}�0�(?CQ��S���!'�Q4+��fs�^�.�\�螑.ϳ�{�o^d)�2�I�Y��l"�}��،_�}�̚��"!�ƱFE�@��e{�a�����3�Q�55���&�.����v�mE�I����������-��Ġ{�)���m���E)�Yf`ʖ@�2�,��r=2�� U��d=��l$GXN:wD��� �'&���;�-����wT�d��A䐃'
�Ɖd1��p��(ɽ���t�yo�Տ���8�v,?J��K�C�]0M���0�P*k[#�!�0&���!��o	���0�,$����3�_��Z�ie�R�k�`�\����ǜ�Y��g^���5��S'=n�SYL���7�@*�]�d�栘A�^���ن�A�����d�C���P��ן�Q�@;	c�3�u����F�h��/���:�yT�mG˚��I	[���>'����t#�)����мf���|ɷ.��'���I�[+�8I�~H#N��jX�ئn�)��Y;��~/K�#�n��%[�*l�*��/?-������C�٪�aГ�g�A�f��H�̪�;�lIs����'ja��b�ҼR��MSdg�B�T�$e��9��w��O��v�����7�]oP��H�;j�=�D��7'U �]�P"��MP��V��R�}��n�M��H�$\�
�Lw_���|0�[/pt�<����ȝS���:�,�2�.���M�6�5�F-�@�VM4�S-гr�.Z53�Qr5����xڜ���A�b����Tر��N��x��.3mS%g��&0�&N����<46��(Ҁa+�ކ���Ӏ���Ք�X�Y��~���fe���~��պ�.i!t�
�����TG�����LF�څʊp��$<�]a�W8'� ��4�f�?Q��:�s�?��]r�T���?�A��0��nޥv��7�ұ/3���4danh�Yt:��(@�:�p�G�O���P��Aؠ,����^�g,�-k����䧗#u0��߾8E>��R�I;%}/z�e�n[h���vOH���ɧX�v[�z��`�Xe�%��	�biv;�.'��_V_��3"��_�A�NS�.��H0��`�b��O�w�o��TJ^~�|cD�NI�7~��Қ�����\��U�e2���������A67��Iҿ��q�pc��9BT'��f)ߐk�B��1��z^
'~����;޺3Cb$	��H/`���o�(C�K�\�F�e�iBF=f`���?���)��3��8�m#���ϋ��0���7L������N������J�̿E�٤����E�f��8�O�/uՋB�b���> �Kx Y����<������g�Y�;��C!yݤ@��.Iu2�L��BO�g�-��B첿I'�V���*OIM2@��Yz�(P���;΄��g�����gu��( ~0�*D��9 �/U�b�L��O񀺾���<M)���!��y�>�C��q��#v�Ҍm��^sS)�5�u"��L�
��Qk�I�dR�x<t�����^j�g[�D��4
3Ff��?��6�!���-�|��A���_���� 7|P&Χ�O���Qey�U�}�˽j��a���������""pQO�1��y�F���O�~��oK�<����Ǡ�Z �?�ے�"�R��Nd��;�'�U&�m��-���G9�#cr_���?Т�h_�-�/����և ���h����/��j���cZS��k���(u���'�$��QOM�3��\�2��x3�kC�Iv{����[��=��*<�����J��#?�0�Ϸ���Z�R�<��X����J�,�}�z����DZ�52�sq��FKJ �nF����������Q���av'۴���|텰�����!��t�Gб��m>6��	~�vb:�����!7�`n��&!S�%���o�ΐ��FqO�T���ՠ����ecZX��;(�i��,���\c�@���O$��U柢�,S_�"F5IF�3#�M$�J�	��00����f��a����ͷ�e���ח����1���G�I��-�
�t�p��;��7<P i���2>���P��c����b��`����Ƙ�C��5'����g�@4��IW\�Wdr{��k^Sl���t��3#���6S���/��<���(�sN�o�pַ�!�[�aL��Nn�F^!�d&�>����Q1��#O���#� Y����I�Cg�Oŭ��j��=�hy4��^���z��ᱴW��H�?`����f�QB���|LBU�Y�X��p.�SG�T�z��w(�UD�a)Sk5���G���}P�wv�xg�������Gϭo弛/grG�Du�x6[���1��Q�ط�<�o}A�Y���<�B�ǌq>W��9��p4xJ�s��w�B�+��[���0ǐ�UIm,#a@vLG�2U@Q7cK$ˆ%df>������H�TBZ�|O�e����X����j����bϣ'3���tzTԕ�?֮h7e�JIW�;{�2 �7�p@�\[�؉��jo;_5w�J��q�<M�u����x�g�+)���6/ƶ]�$�qn����ft�3���S�C�f�揁���yS������!�&���;�s��Y����\VI�8p�ӫ���#��'��Ci��]��m��2��w��Ȩ����X���E��꫔\��UVg��	��Ѱ`��U��zH���������0