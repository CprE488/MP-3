XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6� ؎�c4g�1���
U4{֖��[�\c�� "�ouY+�"	� ��ذ��S@�W�D��:� N5v� ��#���棑������ai�ˈ;B���{�?G�L�(7�4���00��% t��S>�b)E�Hx�-�Gd�&���œn���]bߩ�h,���C �YLp"�c�Nx���?�R��VȲ���`v�"�R���H��5w��슿��y_c+(��}�6I���W������	Kr�����|�r���4n�S�첬�8!��aX�Е��j��u��PL�^��d�������MWFi������!��r�l�7�����RwI�AX~�i땿��ٚ�FC���S,��?;(yoMx*Y��?�I�����wa�K� ގu�_R���%��4҂�;B��F~��a�u�}��$�9�VB���M�YPo�%0w��G+#4}��O�V�n����s��O�}A��.~��'�Cu@d� ���	���E�|I88GU���)��VOL�q�_:A`?{�#�ա��t�`��XNn�2���(��X=��Nc�|�E w?���]�m�ؿ߸��ۉ�+�CU'�p[�#Tuu�������e���u��Y��WŘ��1��Z7y�t�Y0N�l�8��^α�;v`�w�7Ps���ԘO�	~xK��0=�ʾ-��:������W�dx
v��htgNPqW�EX��z��sq%�R���;d���i�"����Ɋ0��j�CC��-g��XlxVHYEB    39de    1170�썻��rۃF�L��H� 6��~������P����������E�h�̰Ltò�����:	xm����"�<3�<�}��9�zۚ��H��5\UڿZ��E������1@�s� �����fB�� S��㳴[O�yĴ�bP��gC/}��]SOp ���?kvP��n�90�Ō���N��j���B ~ڣ��G#��G����v޺��5����ʇ�Qi��KN��íp�A��<F�H��	��Vj�f��g| �4"`ՁEg��������R%�xC���>��Ḵ��j�)4i{�!��F\����밁�S'Î{���eߌ*D�w.Ss�aom��Mj
-):Ѝ�?���8G��t5n!m�:��ۮ��n�xk�E�g�{@���.�T8�b&�i�[�A;�G��~��o�i@=�������آv�������U��c�n~L8��)�(�
��s������b�u�=OIq���#AC	Wv �v�גY�4��S�SQn<�碁�;�X[��EiP
�#'�	MN�{h!��c�m���g��>�tq�b���B�l�5��r:c���5t*,��w0')��u[�,�;�ziU2zL�;��%�ȁP'�W��j���ܩ*n1i�2����zׄcQ0��Ft�։=����G��.j���en�	z�J�V~~#G�be�9(�wґ�}�[;�����}���Q�P-�>��4�U](��)�Mi��s�gD�L�oa�@x1o�Oy���.�~r#͙�wӌ����JM�<Y3'��#L;����b����M^����~0>��r�ѵ��}�,����Z`X����\�(�ʘ3`c�$B�n���u}�#��?�#�U ����PƬ��
,nH�����m�:� �@�A����)�@�wW���OJ_����Ɇv]���&`�7�Z2�+$E�d���5Օ��2�$�d�!�4A�K�3CT$"zO`fg�HcJ�S\�Y�(� ��<�v;H!/L�?P
�l�0�%q�o/ԡFG#��:�Q�P�r�dD�LE���4��.�M�G��,_�/'1uژ
%NF��7�hvFw*��{��q�0c�ѤG�7��%���sR��t�i�͉��[9����BR���ǋDF7mT;?�Z��a)MV�_�e����YQ��������Y��q�̖���֤*6��Lz�YM?5�ۧ��%�@��^�{4sc�0���.J����>��ڶ�-��0�,�ᐕ �������R֬��F��,F%GX��WJ0ͳp=n� �.�{��S����U���EK�t��l�.�����]�d/��TH��X(Z66�{#�%�l�	�:FG������e���I���gt�. �$`���C���w���@���J�����k�\�D�L��ߒ�YGh\Yk�B�}�C�G�;똸��t��ǜp����7��j�pv'�f���	4g�ж?���f5B��6�|f��nj���]��υz����"<�b���Lo]oJ��0�QZ��f��+�Nk|'��wfI|'gH��]q��C�s�SX|%'��>����q;����3�w�g2+Y��7�6i���W>}�G�a��� �ߠ�o��t��~*��&��5Ԃm���x��F�j�9]���_�(�[��19�x�0���v>�RQQ_a�C���F�)2Y��+g�SQ<I�P��\U�OZ}L��9�T��sd�S�:%a��/Mk����:1y3�}c02�H^z�jT��
T�Eǚ%�}���80�{u7E��z����xIR*�����x�Vm��I��;^���uN�:�cH��.,(�w����;��=`)�R���V?o�7���փN��E͒^te���ߺŝ����P����J;��>��W���"Z���|�@��$����Î�����6Nw�E�淞x�)�����7�uݏ��>�(�R��:�i����n8j��{�,��x�����E�5�Kح�h�����hY$���1�cx��:�n��!�zG��1����Т�ATLR#(�t�.�����c�L��WV2>�g�ϵ<�B Ϥ{���^��
�J�p1oR��fఓNʬmŻ�"+O�IY���j$�g�ʩ^�οu}�=kE�5�@��E�yzf�&)�S��߮�7\׏������XhyӢ���j�U?ڨ!m�L8�ݲ�#�{!���|�|z_���(��� ����ͱ
Irv#F���ZQS��\a����E�{�~���H$Ն����=S^vu�Ì;E��@�$���d�h�X�e��LMr���.�72V`�����Y_�SM�A��1�2?3n�n�^�	���ή���]F�(�Q�q���0� ��3��Zzl"���T~�5;o;�����7�NZF�>r7b�y��a�����d��|�8�Y���H�Pbz9;Z?���+-!A�<��h��a� td攡�}I��|S�OѪ�*.�>\�	<\�o����skW�ԩ��{��N�ir�w�E}'�J��P�Jy@1Ƙ7:�Ep�~7����mt?�{��(S�j��|*�W�uo�7�DG�=�##aZ�ĽO1�5k0�L�=�7��5Mo
՟U�U�OR������g���¿;�"�KT��їk�?9�U�A��D��������l~����zoKo S�G%։[ŭ�nv0�^�,�s�5�?*&Z�H/a7+k���Vؘ�̙Ɏ>v��w�Igo@�
F���d��N��+��x�XȄ�v����(�-b�L�6t�������$%�N_�\1%�t��D��� ��֠�P������%B+Yq�h%�N�x�R|n���9q7`�F[��0���� 2�wf)��C�&.JW��	�{��~���?5�̯c�
�Y)�'�cR��S�W������GU*D���]&2��	�����$��	�R�LUp6�T�G,���	��kl��-S5�����@��7�5wc���_��UV��*���B�ȋ�H����Q5ɽ�+y�7ʥ�Ǒ(�?��6�*�yp9b����p�,*�"_�����z��3(��郅�W1s wg�y����R|Tn�R��N+x5`Av���!������2��Rg�d�c%Ar���.��w���K�'�ꕘQ��k��}���.������*oU�����UR�Z�[t�����,e�D��W?�Hc�}���;�Ê){�Fc�Y):ñʪ��f�v�c܉W�����������fa)����"���������_�MC�~u����Rg>X'.~1"\�=�h��[�P�fT�S�����,��:��V0�6���q*=�v�zuy"`��~�	˨��i5�ċ[�e�>��4ċ?��D���DP=�/�֙7ZjHE�~��d��J�1�|M ��+��}�ka�6�������_�hٚ��{�v`��6!�A�;�
���G���m��1�F�g�F��o��\ M-�YTh(�����' Ҥ/��G�3O��Y���v�2v����N;��{C� �@%�x��F��a�[m��:HWVa��6p`���T�D���b} -i2��:I�Z�cn���s$�F�+=��s1|�Z�(�:���cx�x�'�l"�l���>q���zyڌ"1���,~Ŵ����߬��ֆ��ʍU�ZLq2��ϙ�8�,����ٳbiM,er��m���C�k���'��O2�ǵ�qZ`��l'4��|��|�Vy
��df��軦820��-��\�.p)@����
���^��L�=�'j�`M��{�Q�X�u�@\s�T�k�I�;۩.�-c��x�gȏ89L� (����Ǔ�sk�F��>
���U��_�t_
�d�a�?r��`����f��D���f�:Z�j�׭$��ZXKFL�ﰇ��K22�9Nà�����Ks��j��M�X�����c�CIձ��r ]����+yy:��7���R�4���G��d^Zm%�v�I;����կ�����r����tr�G��a��٫׼X��Ԋr���'���d�s��1��G�%��B����\X��K��_/M�`9~��hA��4�hü��X�5�*�R���W_�&��W�j��2���f�U�-�4��d�r&	Ŋ^�[Ra��[Tq�F� p�d%������JU�$;_Y�*Ҿ��\]b/�D�maYG3�)����=<�$N��]����-��G�hT`F������$���힙�"�2�U�;����_�QkEz�EE]T`	K0bbP���q��hP&�a[{���++u$��Mr ����̽��x.q�NՃ0HZ�X�z���XB�gtT�M�r$
Hԣ�wa�^��ز��І�[� ��