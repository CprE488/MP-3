XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ٓ�%V/�U$�~�v0,��9N��u�V# ΰ8����~-����C5{��B.��b��_���K��3hH8a�� Sm a��y�`�M"L��ܑ�_�_ײ3���3R͒3]����J�_���]ez3�i����b\`����ereS����n8�5K��<���`a����%�ih���ҹt�z��KdҎ�=��<�.r0���A�Np��Q�'C��霖S�qf�5�7�m��+�*�+X{(Q����4XWG�+L%bz��=�dO�40_�+���2�κ<.Qb�(`�e��R<�̉Ι�Tɛ�����fS����l���K�+W����NR@��r�
�[�S�v,v�
(��<�LC>�X��*2p��P����=�������Q������	]�s��{�1c�)Y��#�JZ.$[L�R�+�-Z������O��wI�ﯙ��y5��9R`�����x�	"����	�YE�@���<!���)�����d=�Y1%�Е��%�f���13�
���X�j$U��UU���%�ut�\N���^��֐,��P#߯�"�+Z�β!���������aI^a�KaHw�[x+uE|9��x#��Y 0,v	o���JA��T�$R��L	��0
/����&4&��GQ�Ra1<�[�I(a�[�g5�9j��a9W�n�JA0�e�(���'l�]�%��SC��׈���Z���P�7�F�����EA�@�i/TQ.�NxX���xm|/o�,�j�A��XlxVHYEB    1853     810y�^�\��Ҵ㴪�,%��Q?�M*�3�5K���~�hf�K}��֣g,#� ��u=|����X�h�Pxl�:�HQ��^�+=���x�w?D��cȉ��5���-јK�y���#�8A�&��iM�Dh�^���t�z7���r��@�wA�4hk�g�("zܰ�B�l�1Z 0���:�S��4�ۍ��|X7+j)�U#Ro�\�Y�1��E�J���)�X�iϓ�/��g��
)�;�~� >Ɩ$۞�]i�����j��1��
����'K~����N�֊PM⪚5,G[>�.2�����Js6e�e�ٔ�y�!w[ů�{3p�XQI̍�<��T��� �]��A� ��X�ݚt���#�m��0CO:�>� ����6���x���<�M4<°
-%wJ1���+4�q?v8���&�������M���Ln�p�����z�����>���T٘�I�앖��󭳷��Dѳq�|ڬ�ŧ3�϶v}�g�:��ʖ�q���r�|�O.�c��M9ͱ����n��O�"Tq�!M���Y� w�X�{�*O[�Lq`��Nk_ޖ>�@�M�5v,HM�,� 1w�C�ԇ~'h�<���x����kZ���a��@+ t�e���}���<���I�O�x [x{Hߢ��X� �1�.w������ ���9wrOI��$���},�b�����Cэ��#��*2�룎~��f�c��N�굻�δ�$j-�@���Ǡ
ߜr�b �"�0뷀�.s�T#����G��IK���ՌX�;��s!�a;;��@�Hx1�����l*$��nV����a�8�E��e~�D�.KO^K=�&*���ڍg����-P�)�hfrJ�p��{YsP�e�Aq1w���ff��!C-�R��Fa�q����wpN�*N��Ʒ�=��<�,Rl@YL�*�q��9J
��	���݌*k��h�R��x�uK,��@�K&�p'xRX%�]�d<q�+���sv+?���˝,�[�r{ͨsҐ��ha8NH���K��~��%��eay��R�C��B�g��p<?vs�6�|��}��#ʀ���x�}�M|���g�q�<��+K���IB��o3��w�4 ���
x���U��R��,n��[WvV0� [IGo*�K.��
��ޥ�\=�<���;��%f~�[����Xq�j~�����b%M��DI�-G�q.������AZ���:��^��k%_��>�d��q���D�G��:�𶗽��MMZ������;��+r�a�ݝfo&w�]g-�F��zt���]*�!?"�C��/�ʝv>���"�X���V~=/��y{4tϨ݃Rkd�;c~{Q�|�8ĜdkB�V&������.����������dЫ�L�Ú���E����|����;�KPt�	я��=�[���C��z�ې�Y�cF���!'�2�x�vDe�<�t�i!t��@a�Ȥ�l��3��Z�A�V��H&H��Ӫ��Xn���C�,���!���c�]�!�]Ղ�d��������ȍ��4Hz�����¢ܬ��ΉY���&�uJ���l+EI(1�QIf�����c��U����ֈ!�6��|�R�A)a�?��:@��6R$� K�l����9ۼ�T�)��$���ݤY�={��W����-�Y���ϛ�띣|�OZ��\�@ XHg�n/�б޳�A�7��o)������q�3K���vE��jVՁc��:b�y�l���A��MoEŋA7����"[�cT?��n�o�7#.�B�ӭ��\[*�;��2t:٠�ԽQ���L�~�o}�44�n�+��xsf��0�[?���I���X���r| z���m��`U	�T�������cH�sQ.cM��"#F�앖�������o�?�g�9-ɸ�1R�[���d���&�k�}׾�q�u�r.w�M)z����dac����D�2�~~����4��UJ�Ú.�ڍȇ1�9)�Lʛv