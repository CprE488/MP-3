XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���**191Ri��`���p�C�U������P/��B���)^I�@~����NV��˯��_�cG&��
���8A����'�/:&����jT5�~���}�	K>vM��=�?'�ђ�I�BdvUz����a��=��j�J��h�����ب:s� ������җ��᱊Nv��I_�6�*�f��PB��a�J�n��4�����,�fyGS]Q�v�����W�n�?�����'�	��[a���1�fu�߬ʞr�������϶NQpW!�&��/#%�A1Z{�]�Y�sP�N�߃�Q��S���<U� IA��pv��F@,���zO���u��QU���m�L�1^'L�И���!͡�>}T��9a!&6�:�(.��,�,���v�Es��9��G��Wu2�?�s�l��#��Eǧ�?ZvYG�_�X��a���>]�k�A��F�$�2_7޽��/N��~�.p������0`$$�)����-	+x��a Jj�Ķ�s�꽲O��%�ϣs}���b	�㠽�A8
���=��%=�����V=�f�?o'�W��K�&��\���A%��ą���;���%��:ƴzX��4��Q���t�L�H�B�e�`P�r��e[�����o��:����=��6E�AgmN�k0@p�v�`�I���ˎ2��njb&�sF牶�Z'���J����za6*��t����z1�  �2����7�ޑ����XlxVHYEB    2b75     cd0�W?��sh�p!�������:����o�f�o�A��HiM"a5DK�
:$;YA�lE�t��tp|#^f�� 1�reTs��i�5Z����P����<{�X��:2�\\����8��چb>\^�y����`$+N�.h,z�(\���N8g[KQ�HP��L�?�|��"J�'�t��͵`b��.��.��X��� ����>E���X�	oA�ZC��' m�2�	A���,�_�NE�	Q�)d�CF}@��ddQ�Ƨ��H~��M�m����E;B�`,��aT�B����F]L�x3F
B��4ޔ8��ߔx�E��o��6g�CW��'&.��������]�BRGF���k���I[
�H}��m �x_��!���mh�>v�q����ڭ촍2v��,c@��'1��#��m�|Qiޜ6�v��}��r��)k]&�j����J����֑�0��RTb��{�\��� D7�K���Y�AI-��|��W3�;n���Cܫ��Z X�!_ 0=��#Ie�0��=xJv����s����~7$��P�{��|���܁��>�O�J+��i��C�/�O�������Ď����	��J���!vP�\멉�M�/��<N�H�G�B)JlS	�=�YT!��g�~�S�v�$�(P�TUH�����k��f�б��𯘪�puI VU�7��K�|׋�3���m�aA�I[������[�vb7�Q`����b���ʙ�&]�5M�$jZ���{�@ՓYz5�Y
�[4�t�|�����V����lJm�G�xn��H%Vy�C�9�W�Q��0�r(�[��CQ�ܡ�� E)�Tl=*_ɮ�0�>���J������1
���,����u���"\@�>���Ig�[�b��Cn6��@�:��F�=+#s[4u�Ν�Ȼ�SJއ����5%�e�ݪ��B,6�4�t��5���)�f8��Xu�7���H�Ӹg+�||r�@�4�b�/_�n�WKb���Ύ�/��ۏi�y�ܹ�uWÑ�<r�i��JB��k�ު��tӊ)EС��OP�sX��'%Y�x1d�����p}o����@r�W�[˻�۷u�['>37W��fu֥����B�X�Uk�Z�S���b2���k�G����+����J�:	מ�:֊�(�k��!��˅���-V���$����{�fVQM���<28/f�e?��cQ�-��F�"�A5�}6�$�Xl$o��Rr�hJl�>��?]?܀v���lE�ې�sD]O�HW��8�?98��l���#�����q�܌�短�H�y�u�U�j𓿲�
��9�w�6���[�+쉵�*�Qʁ@�S���`�������p���S��w����^1U
�+#*��6��=��`$�O�z�;�����e�޼�\��B�)��-`r�q�������#���h?��i7 
4�k�i@���fS�����
��ì����h��O*�q�h���l�B~��|1�&��w\?�Ɏ%Q'��=J����y���_��`aP�g_�o�O���r�{ჲ�"���i�7�����j�I�ʏ}�h%j����3��O��>|����a�#�F�����z���z��Y��M
1#f�,m��8B~��#�=u�X��}�9sܟ=�6n��U9�ItA���Υ�Ű�gg[Sd���O��t��ԟ_&:Dl��.>�����3~�οV�c�WxK��
i�Fz�;<I
�1/}�z��F/i\��[N;A�p���0�[���5/��i1�8\O�U/��'&����≆K�ذp+ذ0�/q��9�G5�?�0p��+,��'�����
���1�G��#_$ç�x���Q� wP��L2`8�@�P�\�`�D�e���v`b�/&�(E��|�χmj��㳗���Z5���.��=�Gt�r-��?�؎O<w_Q�<�G2�a����=u�\��F��T�A��O��a�~�9�_���7DXe�ʬ��_$d�II�p�z��O�(�[�� 1�z�O�!�X
 �ǅfA�0��?<d��ɀY�*
��;9�|�V�x�)���Z*�ԩ��al$�URK]��4��I�4��Y��Ѕ�:᪲a��1�5c�11��]O;ȓEI'�!�R��Z�|�3X�~��w���A\E� (Nf���ۤ�N1qo;&P}ْD/��G.�$���uMfdqozMwov���(�|<��?&�)
�G�[y<�a�|0
��I�Rt�ª't��u��^S��b&Ow�I�E��0��r���D���C'�n�e����y/�,�u��f��m�W�2oOa�fS�O;��ZY�1��x����Vy�'�i��FK����"/�[�%/��n��ْ\��Lŷ�Š�Meբ�t�2��Z��Y�{W�;S���i��	��3�8;��\|2���AX���W��&M��ݹ�v�|�p�ʛA�!&��K���YdƘ��ٷ#?��$9h�<���A.><�p���P1�������p�o�2nd�k�֋�E�k=��p�dmԝAoH��{��R~��d��@.`2�̟��m�����>�v�h�-��!GF���g^�Q�m��Z8j���34?������Ek��l��]�?���y� �K��oN���W��∆��'����LW��Sт�%�B��s?x��\��r��	%~���=ș��g8rګgX5p�������//���J��]`i��`d��?T%��'�l�H!�VB�� dV�d��{)��eʈ�Sx`9D�w�5ɖ�+{W�SktP��~&��a���|�Ca5S��J�?�o�������ܚjs��(s��i�X:��W�VMvQw T��&pU>E-�S�^�B4 'T�g�����įe�^����K���p�-E�P��\ZpU|�4��GQj�i�ka�Nd׍�Q�'9B�T��S�Q�3*<I_$0�v����:v�6O@H���rVJ��Yϩk�Qg���iq��j��^1~��;�} d�U�<��b��U�sBG�9�t��
��؂�
�7������WB��-d5n:-d�4��/җ�Vxn��ء�1�1�ɋ�U����*[��=�2$�����Ql��z���DՑ-�����>��)Y���TN�H5!{�C'��2 F=�2R�R�v��Pp5�X����