XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����&.u��(��Xu&�������J���}u�c�g��oI�{�v+� �t��{�S<���\�lnH҅q>8�)TW��z �6U��$r����ڢ�b-$�A����e]^�rNi�q�a��PJ�m�I�4 �b��ŉ��N�����ǋ�v�`���3i�)vN&\�.��l�_j�wf�m�Z��#����Dt<��y�0���)�g��2�`��C��ۤ«M`A�G�cf&ܜd���  �0���|�!�8z�8�����2M�V�'Bsk̜[Ff�1�5�e�i>�m���ƴ��|�mĨDӸh�����ms;�d4������j��2ZG�`�m�A(^�tE�I^~��qO�8�$�V��g�KѪ��K�{���Q�zg����h�9Ȳ-���V;*8/�D��P�e�6wa����ղ��X�����:����a��p����B2-jhh���K���x��K$�|�W����kbj�6���!���u��"+ʌE3�<�(�Dޭ��Mr���2Ex����	`bt�hp�|��a5f��~* j���u<�G`GP�	s�R�!�M�������_C�B��XMs�1��a������]ѥ�l)�9/��96�R�:���*lu�� z�t�q��E�=�����	P#�il�@�7Q���鷢��<(�WHW?��>��=��K�|����M�j2����]��#�����*3��v����>b���b�xu���X�P��XlxVHYEB    7265    1660���s��.Vu�bx��Æ�1����R-��J��1���cSV�1b޷9���Ev<� _&$�hL��y���c0W[;��=��A�>��y�Z�j���T��ղ�чI�R�L�Y%�Ǒ����r��a�\������x�G�T�ڰ<=�㠴�L��	�n˳G��b	�@;��ѥ}y�2���FB�9v#jD����t3a��](�
KG�n�͑E���4������
����I��&��H��C���7
�d�k]�ٳ����T+mޞoP��~C��V�A�h��O�GK���XU�䋪�Ĥ��O�W�q˱�h����7�۸&�-P���v��84�vL��2�~Mo��;��~Tx��+��S���_���=��k�����;�l4t3��q��� ������ر�y�qJ��WWF�}X���g�[�R�WeXQW��|�8q�ȍ�t�#��tx��xH�o��_�/�^$�4�0M�2���U]�߯�1	C�s��	��x�A����kBBv��@�5����E����!�|�%|��G#4�M�����LT���d�I��m8K�b�����"}����r���f79�?�8p���t�Bc�.����4��_�����@�3`�;��Eq%�OVY&�/). ��2����z��L�
*�%6d)С�������&�Ą��v��d�[_�����?�diwH���T�a��,���n�Z� ���I��xz��mr�QN�8x�[�Cs�Fٿݒ���ϝd����K���ϣ1!��Vd<^�y�>�ؽ�=_c�dTI#$�q���"P3Z�sR���H�8�� ��[�
�Ms�S�/<����`{�~-e�M�ىx^I�����/5-�8_�q��(Ч$�g$d���۷*�o9������V�=�k#�[��ġ��q{j��� g.�����K�Ec!���a�������
�M�An��4%�=_�h�A���Z��o������q�{�����!�u}vs�h�K�d	�2]��k"�=7&�>)�������u\����f� ��p�rC"(�3����b! U}�{Wiל��#���elg�>���~�N��H�Br]>L8��63F���7��c�2�ii��KW?5�T~D\�"��$�[��ꥱWm<5��)�U��6�Y����p���v�H�Y�,����0� hm��|��v�`@�u� ɺo���I�\���n:R{��)�⣀M����{�K�'5���#�Y��$��e�Ow{�w��U�T'�D�F�Hm�t��J��؆詄�珆�U���ЅIP<�C�p��D��Q�ܗ��������6>��4�VW�^F0�zi*-Ap=Zka�߰r�����v���4(�e�K�;H���D�~�����0�M�q�&L撄�v՞/36�ţD���&��#�쿷!]�����3���֤[R�� }�XDWS`��C�������.�q�3���B+�-�j�ˤ�Yh��ܮX����Px6f��/R�5�Oƅ7�Ç쎃۸!2�˪��S8�-l*�U��<�s�V`H���>�q!\�B���9l!�%���G]��x�D+��Z^�|���,j��6�E�#���qU?���0R�`����&��?��ó.������P�����F{x(�(�چ씡|9�؋�H�k����Ν����eZ�.�M4T�b��I'�%�w�q�C�@�E�*RY�uŻC�s/,x����jJ��{��eP;��������zSȣ
�%�-��z���oh�	a��@dY���lQ�&�d8�8M-.ݖK�I��B{D�H}��c�����L���k�̖Z�+��R1"Ty\�1d>	���u8ڽF�
�0P�k�03=�P�^�7�����"�ff��<Lާ�#|m7���v� �Jo7��!�V�F��ّM� A��]���k����76���!ЮWN�V���k�**������ =����Jv�ۦG9�����W��-��� �K�z�H�%��d�4#�Y�9�0L���g���c�_�o0��T�i7W�mX�H�3��x�xH(�Ub�tJ��
�q����C���&w *��^V9e ���("�`�g'p�q��7�˿��<��gGj�K睛C��DAw蔪iޘS�aV��^�Pa���0Hl�M֦#��P�<����'�Ǔlʟ���1,�ɐxA
}Hw{\�Wsr*���[�L?x]w�fa�!�*r�S\�m�w��_���<�
��ҳ��uѹ�0/�A����^@3�Q�?�w���
A�j����׷��cH3����O�:Ө���εΒ��jiZ7(�Ty��]�+�B��>�����bʐd�;�������oJ�X{�T�F]Y�x�*�1��E��*+?�d��Ŝ�7Sw1�4E��w��K:����.��k��P�m)D�M�C�'WN4�>�綔_ѩ�oX�r$Wv�U_*	`S�d&��ӱ�4� �"𲤤��k�kx�W��%�S	6TȊ����>��,p	�ҙ��EZ�v�&�����I��f^��S�]k���9������:-� )�,�,m1X͢��kmTT��G����|�*	+�ލ֬�݊��Z�����4����B_3oG/�ǭ~O�W�j��kZ�����VVF�^*��#^?����,���:g����e=Dz�i�vG�z�ȝ��f���jPJ�.���F)�$7Lh]Y�}>�Fw��ҹA�;}���Ьt R����+hß�T�9�4�B#ϭ��d{���.�O��
����*$,���Is�/����p�yα�2�D
b'���Ԏ�	v���1/'���1�/[֟�U���PɄ��=� d���������� �	x�i(61F$�ʟ�����"a�ӯqHsi��!���3�)l$C\uf��\��V�#��ޤX=�� �6��-�g9�)*z�����k�٬P������_�#�E��q���1���B�����9�$v�2��h���Zs��_f���Y���t�T�ڌ����Fg�"����3�:c�{q{8��	���y�3\Z�R��^'�g���Ӛ���M����bZi�gsQDG�s�j�í'�hl�F�P/69�q��5�L���t�m��n����]Ҍ���84�[�W��;��rozX�h�`��ċ�ź7q�>�����}%f^��m�\U�A�່oV��]C�L[a�=1�5!��]���oz|�0����p�a�̥�h��s��d�c��3{-p/�(��:X '7�eT�z��WU%6� "t��;�${n�(+�N�B�:�P:u��b={�VdH.~N1���q�ߎ��1���e��FR��z�v���.G7ѭ�1�To
V0iݭ�D�+d����Ż&hU�Y��B6j��L~Ռ��Sm�t�ؗ/�mxd6�^�谈a!2���B�e��%���u�� _aY,���=V*�6�^�Dj����J�V��Mo�u�di}z�8�v#$�<�V>+�����y�V?�w��##Ѓ4�z#�&�5)D��c
o4nM}k �%�'Q}�J�MZb�i������)D����8���I�#	I}���K�cã5��;�4�Q�5zAU��F��ϝ�*������`g"Z��0hS9�a�X��Ӌ��< �^���ѝ��3���+��È;\��Q���"��-���ѫ��������⾐ ʯ��қ�:��Dd��lG�.5�������A	 ��3���ʶ��ɺ�u�� �'��i�)�sePm2ih��
��[��L꾘" �N�b����H��;�(bX�{^�j_���@��O���:j���ټi�z�{��t\@t�I��4ô��I`����D ~䍭6��jG���[��_�;Nu?^����Ӽ�I$-up�*ϝ���b�;�t!CZw�fZŽ�2{$	Ohӑ[�2W2Fц)��R��R�.�d��6�9����2���0Qw>�3>��O��54�P@�j{V�T@���-�B-��8�(LG�`���IZ濤AV5����I��[Y$�%�y);Iz�;I��ަ�v���?{�;,�1�aC%�9�p�G�t4��\q3���ʡ���##Q�ѭ�Ä"B�?p;�]a��ݹμ�X�ž�`~
d�Q�[���@��o"�qWb���/�=	�ja��p����N%d3�?pF^��4-8,Ꮁw�<��Y������eK�S[X���5��2��D�f(�>ˆ	��X���ܭ����P��'���Psf2�c5f��O��hV���Ę��M�fg��	
�wF�S.	���-?���HP������Wz�[��U}������l�Pz�C~"����F�9����p�NRpfL�i�o[�ހNѱ�ed�a�!�<�.�qF���})��ˮ~�N�?.�� �� |8�K�I�в�~sj�w�y~���1"�	"�ϱ�F��{���Yފv:����I�{��W3Exz���;��|b��b����ɔ���)�lp�äoF7lFW��A�r�oA`��E���a��7�ִ�`v�b�B����@Z�n��#��?=s�ѮL;@4�k�5�f���
��!/-�4��O��\��	>{&�#^��H��i!�vf��Y���DE�)Շr� �)�x����}�'Ru˲��>`�r�Q?�m��� zg%X�c㰎�5��j����e��|c8|�/�b�tԀj�?����N�6'��\#U��@�ҧw�-5SaÎndw:�/t���2��e�h��틀�/���v�j��$��`����3�H�v���c�mo�@����M[0"�uMs���7$\��$�zi��5qhO�df��y��,\b�~�jw��c"�~���rJ�����D4- (���]�Ԙ�˼�H�̤]߆a�c4��*v��[�ߒ)�^kx��G���I���,a�:(e7��x�#BI�/P�(ųO�g����>.���5Y�'��#��.HU6��9^Z�4�,|�uLl�D��50�N�<.���ډq[~��V��,��(��5ig���:�iPc�Q]/�:�ĕ��@s�l�e��>z7�0}����[�9�)���v8�Ix܈���rQF�LȌ2v�7r�ؙ`֔E6�oYRFMӧ�8���\
��Z8N	U��Ԇ�S�i�$H�w���T�bЎ���E��(XЇ�NΑ� ?�q�N礨6(��KCɊɚ�a������������-{����$/,u�@`�"�0R�_R���XTƠ~������x�y/�)0[�`Q �pޣ��uvA��B��
!��{�o`������RH��H�1΍������ �:�a`c<��1)<w;ָ��הu]ԧ���i���8(yz#�=��s��
��%��ʌ4gU�̨Xkp]�V��-I-��i�� ��S�o��)4)��]� ћq	�T��� +�$�r��!��%�`Vp���Ñ��yb����c�D�R=PR�������Y�+G;>�$�!g�%$�~UyҾ��6��zx��9�4Ј��&�����%�	�
3��S,�+�{������� qb