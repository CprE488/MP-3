XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����ZNRB	����P2R�z��w�R�0���79ݾx$R�ȃakL�:���hJRJW�?B%pZnj��r�(�J˲�D�k������ra�[�Ʒ(��1�G�!���>�3�p�	,w95n�7w��4�9s�/G8�6�j�`���
˛������
š�;��A�[B�i�*�%�Ǫ���h3�q<ķCs�<.�r � ��2�#*}/t��&���:H�>����45����n��~)�m�S����S�U���<���g��;�	��#S
�Y{����_��E�;�W���Tx�c�-�/�Ν����#��C��Vj�*�P�S �����'ț?���D�5�O��1�D.�1pB����=��3?e�}a�LO�"�����Qj�\�?N|+k��z��φGR���,�x�%>#�~4�Ol��o�Ւ�p�yg�Il�g�/Q��Oj�I��9�����G t�(���`���޹G��@'���'�LI�)	~�|�҆K��J�_C� �q�xE!�"��C����1�֬�~��i��k5�,���K�s�y�|������>�ff�^[�V�d�>��<܀{�讇-C2U[��
l"�T��4 ���A��vܖ�,�O�O���;�h��H:#�Ԋ��k�2�w�)����d�5�?Z���oˆ�ߊ�X�3uD�*��ͫ���*_�d�C�{�n`x���EZcf�@IA��(�)7����$��8-{�`l�0�)5Ѵ ���>�A��XlxVHYEB    1421     7a0���p�9��+(�Ͱ?��h���}ju�Ӽ��n�ǻ�R	��9���Pň�-�ʾɆM��@ʼ����m��e?�lPIZ�c���=����J��̮|��_u�+l�Z���������!�����8.��t�m��>4
09�lu�����󅬤vkH����Gp�˾�t��W��H
��Gnϛ���f��U*ی*��e8��
j��sP�f�Z󎶶�,���;	�K��Zg=�hdl%�#>��|����8�f��ꓑ��HE^��WQ�M`���b�4;���VG˼��x�'(�x��M^�\�eR�C�n���`��K��[G��~7���ؘ�;��;��`��ج����|�����D:h6�c�P�K��1iP��+�y�`�XbH���.���~�0ܔt���;�ݽvz߂�B�h� }'Z�$V"Mp�)@��+�}a���˓�R�pH��k���%��cz:���DW�t6"�(�+z|�����8�4^óD�:�ұ���>���1(}�%8D�[J�=�P���_O�2��<��D�� �KV�[��4v7?-�����H ��\�[q]$����U8q�\MS��)�t��˳w>����F�_{"�o���J{�J+U�Ȼ�����^Q�G�C���1D�v7qed^�dʐy��'܅��#��+�V�Z����f$|.o� 1��L�0��#[�Q�T;N�����p$�cTu�v�g�\����.�z6��]b�([HOaI��?9�p"�d�u7������B@��֥�o[ӑ���*ʄ__o���|.�?^}Ǆi� � uԴ����ػ?����
��w��J���t:i�r_� H��X�,�=�F�TJ�8ы��"�,|M�Dm7ʌ�7��3��Yw���+O7�h��w� d�W��a��{�'�Gk��e����S��Ai�p 7��4�ޅ<��'6�vp�7@ _�]��l�GW�j���#���Hȡy4�{������4$_l���m��1V��6N��	~.,�x�����_�9Z	1�e�CAIН#�館�r,/p:����X�E'8���hjG��	�9�z]���h��5]�2�$0P>M�n�^w�0H�;���yrO���^ם)�h5��%y�2��@t��0cQ��`�����hr#�zuH��g���Rmyx������L��B�Ⱦ�su�MKD���^	!��i���am[�o�n���������A^̠Y�GJm<�g�`�5n�@8�\�� ���X=��t��Z`�n�"�Z�m�j5Ǜ�O2x?��#�$�s����,/��L�y%�r���|�:N!�ϟ$�5�[��Ig�&v����E)X%��6����پ���ur��������e!G�}��`g�m��C⠧y6H~{4 �m=�֫����5�*��*#�U������@���ھ�[��nnF]��T˨����a��Z�j~����I�������7�ė�h��C���1Uz�1W���� �u�(7�C������<�RME���y4B6z�������1�:)Օa�F���`�N�a%��I�t�y��/'����������&Q�+���4�'���
΂���&�ޢ-��c�G�^�B�4ە{5A)��Е*�C�/�/qX��\K�?]`V�8�AՋ��ɧ�[y�q�UP��V�jz��X��S�9�M������L�|�2<|~��ݨ�st�L�_'�,��0��SǍ�[F�\a��g�zC���APV�3�H`���}%�j�f�Up�(v��>�tbuJ<sW�S�b�1i�:���!�(Q��g
lC�&�Ֆ�Y\�#UY#ɉ�'�2��z�ޝ��v͙!J�q�z��I-O�֠�9 ��
9<e��4&A[��K���͙q A>A���EDo0\1����5$�z�͐�~��vN7ב