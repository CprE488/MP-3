XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���T��x�q�?��#M�;����Ecl�C���k�*9�ٗ��gj�msҦJ|?�f8:�.n �2C�,]���(	�����e����g݉��zjs�y�$n���5^;���x�_4����V�1�����)q�x��}/�p��������|�B�i*U�G��+�ν>��G�(@���U�"���*��o��̦�]0}n��G��v�+���:��6�)�*���u�g޲c j1+U��R7���On+���6O����P��p�nJ��<Ia2��A6��
h�9#H��h�)��̄b�'X��fWu����T?��f1D��	�W��AM���ບ1�dmS��Eˠ*���u��R�d�x�;t7"ڗ��5t�]C�JF����֩`�B	?�b`��V�|`�Ի�ط��j�\"@N�}1�	�#Wč7����+$z���fs�����t��G��m�I�m���=���l��O�8;�/��<z"�DH�+��|ۛ2�
��V��R�8����ic��Y},����0���#(��/�оi"w��8j�p���,,sG�maËcZ���@S����vC���Ӟ�T���C2��I"!U*�\f�rB���V�?���]0�ױG͓�y��d����|�p1r;�H���D
S�kRQRd��Ѡ�/�����+8&\�,�c�k����)`~�m�'�Z�� n�V��uQ�à\N?�^#�{�� ��fG�$޹��a���D!��Ԃhm(�XlxVHYEB    fa00    26e0��Y?ϕ�{�_e�]�-��]ht��Ƀ�D�]n����	1ftyi�0{�ȍ��;!@�j��x�����eCe���I&C����v�I�ؗ���L�%\�;�Zt<F��g-�:f�.gȕ+���xF�1ԛ�X���\`������Ȭ"8׍�$�β���0�$l�]������a�]l{���n�.h��)V��(X|;�9	�,�Co
%wb�G��]x�V�.)?#�O��GW{�-�ܡq9P��x]Yw�Ѕ��f}����l��P�Q&���x+�nq�kJ�ZNGn���4č	�_�/��V�85x��e8n�!O*:��m��a�!���D��W�B��i�O��=&d��|�DԬ���f�7~@����XNM����倆(:i��=	`VC&|�U�����l�lF�v�s���^��Ow�D�\u���Ɲ�wg�q𖱓r �*���[4��D�6��Ҟܽ�62�G	;SVY�AT:�ZDV�%|�.��k�9Ny���w�?�0Q�o!�ۅ��n��9z�	)�Ƃ_�=k��.��F)����\j��íLO��#��9�!=z$Ȼ$U�І��A,a�M�ٍ���w"vJ����Ő����a�,��7�ftşk���g���;�r�T�w~B���&�7z�ѿA�ڂ/�����kP�$��9����?�k�A�A���!�h��A55�v����~NokM�Ee��PB`r".M\e�2��p�_>i�NA�jxV2ه��<߿�d�mC��y���:��llo��n��x�I���M���vq*r:�.��^��II�N�����s��?ķq�.��,r�/�BBA
��$��f�7�՗�C��p$Ӕ���p:h����Xd`~>����r3�M��F{X��Ћ���m��B�\�:��HP+��0՘6����	����T�	�E�i��4�&cB�@k��VD�cf�v= ;s�TMשkR���ȱ�O`�%+����f������|?�_i~�,�#�o��O��ˆ��|zYB.r�ث%�Z�tec/I�R�Rad\G�C���I�"7t�:�O������r�Q�t��+]G_�R�˦��N��Jd��ް/?��Z�{$�l�M~��L�D0	���B��1^\���0ҋ|4E��4��+)*xtە~+�ZߢW����?)Ν>e�@9l`��kZX'	"mCM6"`nճ��n�hٙK��_�`X����U�,��x�UH"�b�q]x �38�.�h���r�����gQ��d���S���o�g�= 0'ҿ�qOd\;�r:������q�?;M*�t��~r>���	/-D�W/n�z��W�u9�t��YfHUR��`Ƥ;��ۯ*�y�������S�|�P�����=�U��:	����d h�K�j��;:]+�ם�_zr�����Ek�VC����;/5:���� $J^����Pq�:˶)�'ISA�c�a���&�^�H��w,���Wl8k5��8��Dx�~��^��,]?`Sg�*v���|�ݣ�m��;"�'4^ݸ_\��5���cb�\�ؑ���-@Rʂ��*pT�yx��W��k;w@����)k���}�R��	�ݮz�W*0΢Q?R����K��*⌮��3Sԫ�����.�Rgႍ]���_��{�OsmM^)N��?q�As�5��T�5��rvA5�ANr*���r���rݐ*v�C�~k���~݋ŝ�Y#��aw߮
��DMaz,�3C5.��%�#�h!}*q1�n�0�
��51!��>�;�N�{Za�-��l|�_\���X�Q�|äi�p����BK��	
�F�l�u�b���E<Y�-	�Ge����_J�و����ɐ&�A��|[7B�D�U��|,�T	/�#��ż�=�|�9��͎&�]��_h������k�"9�+N�g��v��?��wd�*�v�x$y`�м?��u��/��Y�f�rC0"p�n��O��U�;��<�H�ڻOy�ċ��Z����
��^�<P��ګ���\]'^:��U���B��D��I1y2O�W���Ȍ�I�(�|p���$p��N9=�,��/�Q��B$�Q���
ʬ���:q �~·/�d�wm8S	s�s4��23�u.	 �Sc��#���!�;��#�r@W�N�c��e�.���@U[���Aڞa���� kCo�Q�dsW`�!�����}<��9�-G�4"F����V̼��܆�N��fS�6>�q�خڹ�-��)'�M�L����tf�f�]�UB~���n����p����N��c/j��m�ۘr+���Uz��g��Y�	��aR�yw��7�#����cEo�w��M!����G����q�i�@$�y���a��k����R`G^�b���?��n�9.�1*?���<e�z8������#;��H�'�xF��IC��x����,�B��哻��(Ȃ��3k�-a������q@���U4�@�U�E@ZLL���u�[&-,Z�/)��Sq�$ ��R�k_����o��"�TF�,eF�+��WrUp�mY�':�ȝ�V�~Q�b��
���0�TLE`�s�ۀI]���8T�Ă�&�P�j�;�N˿�x�:YD9�դ�a�������I��p�D�)p+�K�?=�(y�5}���MF2/m� �7�V�L�Ѧ#g�uv0�$Ɩ���$���h�P*)���d���.3��C]���!Fwǅ7����T�,R�C�� ��"ڦ�P���""��A*�r�����柃7���zm���5z�����&�ҤS*TR��2��8�`��U?�"��@Pi�<v�Ε]Z~_p��ݨ�P�#��C��*�K�wеr+#���k�QM(���~f�6Z�w7��Y�]��E��JY�f�o���H�.Pӆjv��{)A�E�3�x KF�2^A���Ÿ]���
�G�D���E!^��{'����& ��^�p��!�>��/w��.j�8�Y�2<�؎�$��e�H xt��}�̕}�c��0M#g���.r�.RT���`�W\\�������E0����uOq�������md+�3u��#�n��|�S ��\uBA?)FѤEܠ_\:<a?6(�?�����I��^]� ���_���:N����4�+b��8��p�=�:����A?���J��k
�v�� gCb�����4�Yߐ����]���@�G#cI�<�~�<�y3ˊ���z̊a�[��|��rE�qA�R�N���M���Hǚ�Q/փ��&Q�*5V�} ��f;G*��y!���[�?����������I��e���u��5�����4������[�ӑ�`fV�8P	&���Py�������s�2�%)�d���T�Z��P* �jd}�SJ �P�6D�|+͈^���ɏp�r��� ׹ͬ7�
ْ�$��'r,Le4����pj�����V����Ky�l�ngJ(�»�2�p��-K�~`������j��g�C����̝��p�x�࿈��Sg}l���ȗq���hN�{9�7�FX�����2�a=���C�����-�y��UN���|�Q�Q~����E��nٶK�A-�� (�g?��OT{=���`VLO���aG4o�@e(�Vέ�|�����,�a��X�y�G��)`�B���]{j|k����d7b�gD�W��f&��C�4���E���v+��5�O�'S��<�N�A�US_����%���y����rvp���R\�$E����~'�c@Ϻ
��õ��U�����V6�Z�Y�4o��Fd(Hm�e�I�>u��Ҥ�@,�`��m��5@Q���{�0�Jq4�55=��@]�]G�I�̀u���`R풕w)5��=$uB����H)���:%��1����2�LY�ۅ�/���M,����UCN�0���9�2��0��GV��_�@9�ܞLh^0�m@�F}=�(�`j��*��-C����eI�^)�L�{�$�:/�D�q�&�`Y����?o��T�t��*r ?ʺb{��1����*9����s�A�*̖�H������ H+� x�cD��c�Iw��m#�#��@�^��hV8�Y�D���:ER(���'��y��RϏ�'��قxA�%�=V��z�������zd~n$���?��䡸�ѐv���<��|��t�g�d�%</�C|*O���C��I�K�,w�K�7��\��_�?��}���� <A��/�:5iˍ?\r���%"I��X��"��S�#^��\�j�jD.X�C��4��ok5�}L_h��I��a<���I���O2=��-kE`7������С��a�Ȝ~�V7��5��2Q��h�u�C�I'+95і$VԔ�l76ה�u�i�.�uP㈓spJ�ěg��z�2��~�����6���.AսB�!�2�]�Y�]te<�v��3Z)E��@��'�ɒ� �p������&�Y��oc�� 1g1��t����C�,�5Hӻ�&�^�(�[r"���eY���m�����ȵ����?����jG�,�	�ut��x��q�R���u���Oo5��`p���`�6Z�ԗʁy�l�������,���ga(��5�ܕS
Ä����`�l(��� v!a	��k�DF���oFw����#!H����'�W�
t���F�/�9q�?��d����ɽy��k>@���>ʱ��+&`�jf�j���q+��ಕ+\�ˤg��������M�rU$e3��v	�{E���w^4#�N�%)x���¨#&�R��ΰu0e��L��rե�
�6�F�~�V�5��!����߲�C@i���^c�&mw���M�2*��(���%��^�Č�2���L$��-E1���5T�u@�4�v}�	@
�`E
���)y@)����=��F(�s{�"�����Λ70���x_;��;�c��gQu�]�iGm�7��<;m|�堗9���]�4�NYj��pK�:�^�}�6+p����R�q9YLuT��yI7_��y�C��xf��rc��� m#U��7ׯK�g�[�@�P�����M~P�k
C_^e�;s�:�I����������>���)��:��H�n74q@���9��DXR�૎f
�4�F�u��1�ϳ3���7���8��/j�h-<�OI�&y��K:�N�0�MϏ��ƍ�\XXA������+��Mj�݊���JiΜ�t��[*���q���lHJD@~P����H%��as�;y��<>��9�<7xvf���Pa���/\��j}ԩ��sy���L�ɕ؏��#zH���ε�] �J�,o����%��O�KF<�&��v��G�7��3�˪�M�Y�rS)�!t�
\?�j�끜�������(���`d��{��Z��������O�wy�f:�g}zn
��&T�sk��~*,t�I!p���>��I��Ƣ=yd���� 0���S� A)஺�x�n�X����M�d����9Ђ���V���͆E�l���̍�M��UҶA�l�B��Y%ȷ��_��Ni�[�iU�Ҍ�
B�����P{� >Q�6�/�qn!XVA�f�A
1r+U3 �AN��K�����@�E���*׸&<st�l�h7T�&j�R�/8����S`]:����);x����Cj�Q\��qM�7�U�J��a'�E�4�N��:������@̰xq2(}C�r�m�N��@��9|��)���{V<�s���|�	M�a�~BȡpD���֦2���+4	�f�?@�B�րf�-��.�Q'8�x[��2�5�Y9� :�-=�r�d�ݶ�`�k��g� �}�]�F!�r/8�ff��p{�Tp���2G���iU	�g�.�o��l��!�Q
��P�
��Z�&@�Brđ�,�.�N����,l/���NY����;vU���Zn�N��5e�B~,�/U���yֿ�lv���:r�
�p=j�3����k�c��F�S#sca���b�[ς1�XY��k���u�5*�����%.7|��ꇠCG��4����=��;�Ui����2�����~�RK���Zf�j��P�Z�)>�f���/H�_�
���|BM�o��	��P�̚:9�#R ����{�l��ߞ��L ��/�vr=�:�1�u1^OQȳD��4���v�6���|�~�)��JRhς������֓�/Fz�r�a:#l��1�(�B�����u��h����97�sG	���G�x�$�E��b8<�*���rT�.F�"���>�`;��}:Ö���
���'��9QA[�ϛc��j�V���{ r���b<H�6+h�퀍��Bg���S걯xc�=��A�c�q��8��QF��,��:Ն�<H8ޅTvO���`:i(;'���n3�,�~p	|B��Bp��y~��6o�Uu&*ђ^�ڔw ���vh �e������i�i�Ҭ�����LX �-�wej���ڋ�n�b������>�q{D�vu��Q�v(��f۹R��bDH��'��p~�sf�s�]�>Nn�<%^�Y�t16+�$���e'�v���fS���0HsP?Sp.�]*������^�u�Y��'�v 3��	%�2�X�3�/%F��|�� ��>�I>
4��Q��xӹR�5�+~X�T�/�Dqʸ��պ�^yu�.�n�L�0��ۧ�>���B�6���{	��1��ʩ.|�ib���d���9iS�ί��_m�d<X�Gu3����T����(4�ݘ������c���R�J?�Qm�RX���GEĘ�qF��q�)�')Ef;��ޥj�b�W�x��W��H���}���C��ͤ4��_�]>^|{�Ș��]�¿�'P�+9ۻ7VS��Fvi��� ���=�fO��5�������[J������|���{)YG�H _f����%��t�S�f�e,���y�[8>�=�	Z/�����:���T3�$G���+�z4�7tQo�D�+i�]��?6G���{�4�Y�BИdzfQ���"%�*��0���u�F�G�D���NK�K���Ͷ�J��`{���ǝ��sa����k7�;b�%j��ѝ-���븄��l\����������j�h�ˬ��b `���e�] 
�� �
LHTӋ��v@� Q�Ȧ���6Ym�nP�#��Bܺ�%뫭���TAl�S�]�&Y�Ǳ�	�%�4��<Ό8[Q�"�(��
g�c+�y���Ҧ����`)���/+fκCz~��2��fM#+P��F�,�a%����㷯aF��nZl���A
�0�i䊂�CI�����[|*q�j�B�7��*E7��z�A�Ln0u�yXפf~? �%��G���`v��#!	�����HΗ�������_ 3mq�I�u�����ҥ��al�B���TB�sFye�(�����,+� �
�8f,����w�!v���W����U� Ou��z�,�� �<�8��o�̠�K0!��
,
�TI��G�QD�t��b�.�C�6B}��Z�N.�w��(#u�#��9�6�T22ƣ�e|1��d��N����P�wڟ�d�b;��q^�7h�����LDg�O�:�LO]�����K%3���e�-�)��F��n;��̸}�䦎`���v�^.P�����8�d��'=��N��+�X����;S+A���dm{+�%J� {j�0���y��y��[��(,�t�g�%(�I^��s�����#���̆ȪӠ���߼̃m�V�a�Mq@��-�����ƣ��nspϳhj�P�%�(�
OJh;�t?���-�!T��4֤F��7���׵�<D�`�w�G.O�za�������*kE��]���#z[�wzTT©y�u���W8�:�̐���	B���b>������䗀�� ��Y�;w�h)��:�zԠR�z\�ǋ�����>��;[���k��i��'Cr�g��{��(>�Z��w��>>��
��.�-	;�鵏���<�ByI;0@�g�f�3��~�<#��pNMR�c�,߁�RH��5���/��v�����0e����&Bu͙3��vg$>&�-G5_��X[f��п\
b<�]�g���s}���AowQ��T�E<�+'�]�nz�x��9��� �:��v���n�J���6�z/�����Rg/e��Y�G����ќ��]r����{8G6:�ZK�=�'�I��j�m	,̨���a¶VV<<����?�0��/��p;� �?��+E�"�J|�zX?1W�&�%��	ƻڛmw"'����NS�;P ���X��WԼ�;G���}7�V.h>�� B�Vv��g���|ݑ"G��JZ�]23��tȵ�gq�f�\�F]�VJd���Ӝ�%����82Gu��]q�^bs�z� 98b����z�6auNX�};p+�%�[�'����� �^��{��I����G�{�TU�������i���l����H¡,�QR��������\f���=�T��^�\��Gc�����)�8����}�ؾ�[�\�0&��H�(O�>�Kk �[�g�E3T�b���D����C��D������"��^�h�44g�d�
]��܎�Ϭ{@C\�������]�Q�u�v�G�i�lt�Z���C?��1�`%
�׸������(	؟8�e��Hބ3��GdbF�C��.�|7�.��ԩ!����h��-��B��zU������@�����T��5-������?7��$���&�������%�Iz֭Ԟ,5ĉ/�c�b	@�	����SZy2%Е:���5ҷ����OB�{`�^@���
��~*�Ox�6|�Ln�4Fy����C�Y�,�~1M�>���gp�F�Lg�)�l�U�;���b�^جvɝ��E�m�3���/�{����o"���V�M���Z��#�_��������4��,���rE�ǟ�P`I�s��'����g߭K�%��0~�kn�=�W'ջ���U���$=��-���[�ȵ0S(���^�E��b7� ��|a����0u8<H�g�-�ڏ���ؖ!֙<��ҩB��)�f_Q���pD���
�j\��0�f�y��9��\�����u��pc��� )y�h�,������"U� {���8�Blkkd[pd:��e�r����m���BO/K�qT6yd=S�T�H vS��Й��h�S#�/�{(Y����*�AC�/U$�ۥ��̫G����YCY|���G��׋��H��'ʆ�f����m�<���E)�	�_f1����7<�/SxlR�KW�F��ǔ'���|�?�yZ`��z6_�����?a�c��v`)m��.��sJGP��}��hh�(
4i�'��ר�hn�=�������zn�zJT.���m'Wη��ٕ<��Ŭ�pv([�Ğ����ͳ� Yl�:����	d�3��t����ۀh���Y� 9��1AW%n!�Y!�,pc�H�����A0v�<�k
��-����F!���^#�b�)�Z7���x�X�FQ�x�gS_��� ���[u�xz� |�9SmV.[e�ޤ �S{`�S���W����*@nR�^a���u�l֩}�J~ӥ��� �Nn��**��E��+tCմ�Y��a��0��n0��}`_D|�]�%#�?�z򟤩A��AH�Hm2���϶��`�$:�@��S�A�����__�_�&�B�@��1�.Xۖe�4XlxVHYEB    7d55    1450 �@���y̗y���)���Zs�VxQ���$�Hq��o�C�)��D�q��Q��0w�Ϟ˛�}LJcg
U��
�m������U�Q&].��#G��m.� _�@Q����DS��e= �6-6�ώ�)k�Oed�
�V5C�M��h�79U3I�6꠺�I���yp�'��f]�x�D$|���5+����� 'L3�4�/���]y�,)��x��'ةg�e��{<�IEo"�~">E���|>�AA�E�'sV>s&8#����#�2R~�l���lө<3�N�-/����L����;$��mp^�GW4��Z�� 4����Bm�֖��F,;�j�+���t�H|���-	 X���`җ�rJR��J�ԮC��|�����# ����b��x���}v+2�	�*ͪD�A�ˬpa(���0-�iǦ�\�6�4Kn|�J(w�!�G�@o5Ǎ	p�Di �nޥ�Goj�0b��᳥#��U�|dDj
��8��C�r��`���(*���"{Q���3��<rO���V�^cR��!��Mx}�Y��dPL�m#��f�i��M-��Αb�Jg��8�,mL��7�Cĳǟܬd��@�Z^��0���!8;�l�KPzr]I�eB��G,������2yҙ��	H��e�.a�q{e9�W�>jO������#7V�@�Y�̛�|���(,��&��^�5����u*n��!{dP�G���4(G)$�F����E�m��5H���@�N�XR;�������&��}}��]�]BOD���'��]G_��������3��?�a4v�������HLe�b�� �7G�jdA�#��[E����g�D�Y.��{����3�I���9<5�f�D�GCq�L"˻O��g���Ӫjun�t�������B �3��%�?)����ݽ~��T�b4`y�yȥ��fs|@�W��A�l�e'�`5
��,�#E�M�}��=ldV#LR�T�Y�&���Ã`���\�	�*�s���,e�0!Ib���#qa�Z��tG��g���h���^j�V�W��< ��c�)sͿ r��^T�׷W�ϑO��Q(i�N�z�������'YS�½w	7��q��A*-'���9F�Ƀ�7E%�`�dJ3ˡ�^�H�k��o���Qe�����5��Teq��v�+�Z��q�4r�?��?m��n�#�����-�]�4ߑPM�l0|Xg�`�ʄz�\�%E���1{
8�^)9it�l����}F��0�G�F��~��FV�]�M؏�OG1In^>�R���$�����d_�[G���7��$#7C�R <��������14��,�˩����UeV��v�}E����^K�}9�-�}.�%����p*E#�U�=۾Z�L�VRD�h��ݕe�:�જ�P���i�����T���m���k����� �7����E:�� ��l��N$+Ki�V�/.��~���,*�~\H�^����COy�$�fB��8dITj�&��Ef�0>�zy9	z���۶� ��+�
4��,��=Fa�}�3by����$�6���yH;��X�6���<M�Z�I&�Y7FƖ'�� .�ohCb���!���w�UB_��i`޾��QzkL'�IZz������x@뗐t�� ���Kg��$O���R��F������nlaqs�i��8�d���I��_���9.`�0��n��'�1�1�Jz�j���PF��mQE'p���q�S��S�[E�ETo}�KiC�@Ex���BM�|ˊ��sϞ�О#��BG��T��u��%w:��6�ܭ"jD\-�k�EIir�8��9��sű�:K�gβ9�#�}7kjso�,�5���D�k+8�|�k�:�Q����Iu��p~Z[+�T���g%�`E�	ITt�Vl,zs����¦��7<F]($��W�)�0���-�V!��Fq��X_��7��F������ڞWU`�'0K)s�*fq,>ɠ~p����~��v[3�xK[�8���x�= ���H]0�Agxx!oՍ.?M�t���ї�9H��I�|?l��lH�� �@�2(�86�("Wu�z����o2���)XA��1�?=�o�q%\�b�iT���V�"����;��(5����g��ðҺxr��7[�S)@s�j��D�7�D\�N
��Oo�S���
E�V�^�x�u1	�N��s�r��ZHa�)��;m��(`qtm|���Z�%��6�+�W��3���a�rD"�?��F��ȥܯ����ޭ���r؊� �D��(��^ZʙX�t��eS�j��ai �Pp�͆w.�9�:!�(/{θ���v �[�������R�I�*w��ak�F�����?VW�����	^���E� � ����5|.=��Ӱ��L%��j�J���ҁ��²�<������2�Im:#����qU�J�s�b��অ�m"x�pvu��y���C�m)�$b<ƞ���Pp�?A� �@c�ou"{��SmYb� �N�-��b�e��O:�,N�-馎mӮ򾖵u�F��5�n�.3������y�(n�
�~��|-�)ˈ����j�@�����W���n$�G�1����׬Q��h��^^�Ff��̲>�A���r<S����jl�^[.�Ur�>(� (f�@�٬%^�hXh,&4��m�d�l�t\����>M!l����4|�����+���H�R߄�U^Pm�E�àD�q�N�wN�05��Ou�r״~����
{��Om��RUY2V���{�0<yjzX���"���Cϝ�=M��	R���M��JLb��;ee����+e���s~��s��!�ʆ0�C:RX�Yr�Jd��%t@"�B�X�=�[�d[U�W�bܩ3��br�����������ӜS	cĴc�=�C������^g��]��$�&�mĜ.��ȥ6�9Xuc/>*;w��H���y]"g(�H�~��hk"����M��)Ag�ylb�+�*��wt�C����D�s{�,�j��[(�k���8�|�eWfM�P.Y#�(�#�^OSf����"�X}��|z�/
��ش )KR�	D1��#$�[�,�����
�@���Ck�^x)�~����4AvK8�Ȯ+�(`T8K��Җ�m�+Y)�z�oP�fH���Z��D��_���B���7JO�<k��Y��<t-�)��R�޺��3��5~����a���ʆfq*�s ��R4��jp�BI���8�.�H�R[b����h��9��Y*��t�;D��� l�}�S@��D1����)A������v����	�m*�JB�4o�Ź��e
�T��x�E��"Sf�+ћ(g�Q�Aø��8�B:p������I8���v��f���-�k�n�I���4�Ӑy��)}������*�r=�5��ӂրa0h^�8� ���%3�+eα���1j��[���W,� �f��d���!ͥUֆ��$t�@���u��dM���2�Ir<�V���
�_ռ-��p����9�5�l!�*�va���mS;ȑZ�8ʯe�~l��SRG{9�+n�FV�2�-��zb���S\���#g��ׄ�;
��vr����5[��}�Vbf���TF
д��N3�'H�y@�yg��pG�ϯv*ۏe:�����U�_��h��W?ǈ�k!��)�Rb�D۷�%���־�`�(�y&͓$�!.��/�Y�IT��zI��x��MgT�F���m�j������]�5�����f���7����#��gSH���;�m@��U/�seē4�\ah����\�s�Z�jd+B�%60�RUy[����Q���H�x�\�W��`wm�U���A+3� �QM���L��у�O��&����g����Y�T���� �P��r��>Y>'���?���e��N>���)+T�Z|q#3�6I�	(U����bA�=P1i�������8߶Jz�p$>�����k���s�����=i�>�\����4?�}���[I�L�z3����c%�_��~�WF&��R�}?��uyx��]�FQq�ѯ}��<�p���P#ŉģ/�e�Ѿ�'3�À�E�@���b�I%�o�� �/���AЧЉ���v�r�Fyϭ�Za9��Z�d�7����}7ǧ^w.>A5W��+�8S�c���2w���+���U�[q|Wo,�R��q r�)"/�s��f�d�o�?�Gc���"�Q���I;_^�0I�U�(���`6��q���E��?��x@�Z[�:D9�
A���m�B��	0ldd��x�xd�v.F�Qe�=}�r(�c<�΃jVȓ�����gZa���zݗc�LD��ʥ����^LX��g��]l0m��g]V�D�x"AS��gXF�Rn�!1�]c�����e濻�N��cs�B}��MD�9a&�s�Z�̉LMȾ��7p���:��  �f.2��S����oh�v^)A��v��b�ȓz�l�_�K�kh�`��Ϸ���	px������yL�Tc�l~^��M-�n�Gʻ�n���I��U����&��
q�ǣ��,�V9����0W[�*�����>�o||jM�'jHlp��Q?���.�܋(��ߝ����7��&�Z(l�n�SD��;c>,��s5��N�U�҉��F�I!�޺i��?��Yx_r�pVŞ����K+[Y7w�18���lߙGWp^!"�c	<�m��� ���7�i�Q�M���<�T� �b�W��|ʡ�nkIIv8�r\�}#�JI0:�~i.XP$�q�͒Z�VSe��d����#d����7p{\�!{��W���9q. �"���h��זw)�˾�x Bm�JQp�$Ј�+���� K,�E�ԫ`) ��� D�9?���y�[��̍���f�>�vhu����/u��pV�z�Q��Pψp;x�/���?H�-��W[���y�6��_��^yCC�xe���}��s��4��������v�p�<ƥ�P�By��z8�*4�V�� ���������h��}��O?�\�d�atn��0R%��