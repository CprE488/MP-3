XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���i�@���Z̚��ښ���kqo���U����FUS`���ll�{�sz4����W�;"���࿜���5K�9�1ͳ��Sö,�NN��#a���|���Պ��^W�ǚ@p�Ѽ�+y,|�d^�t`"x4���	����N�
Ue�CRbH+O|t�)�"���D;��2�F�&b	��S�$����`;��x$r��
��/���\�(�Ln�9	�����Z��@�������u�iP	�Iɖ-Le��g����>D� �+BTV6�M�u�C&�;��m*���b��w3�����I}z�>�ƝI1q�EõPP��x-��Jq�熙���3R/��ɼ�e���QM���R��� ywA>ښ��"�b�|��V� f������x��7������� �v��0�^ы8��L�p��)�p�����Fm�7�=�۬E�aӎ�6�[�JY��g
N��D5j,�K܌X�Eޅ7�s��<���kmHZfҐ�8�pqmZ��R�z��=���H�&n�4H�	��� 	d�@�	Kߗ����iX/������_`ov�	^��@�:��G`c-v1.GB�� �æ�oE6���OZ:���b�7_![��6��fdP��f���(��L�����Qy$���p��f+��Ʀ􏁲�m�xz/
&#��C:�s_�u`J��]5�l�G8{�����N<��kT�g�o��o�vڭ^e�7Yّ1��^D;+�5\ʁ�A�������{��`�񙥅u6/XlxVHYEB    95d3    18d0�I'�a0`�?����H2��Wr�+x�Z>3N7�la�A]�y���ZnyX$L���G�AuZgӰ2r��2-�۰���wY����O�2�nvRւ{���0S����_��,�� '���.�Ч
q���AίդW'`5X)dNeQ�0m\�D$���Nnk�^pϪ��',UUr��."�V�f:"1�'.�9���X��M:�5�=a����[� YeV�r7A�-�h�D�S�>q��6��8h��Ѷn�
A0���ZEm�3�k%)|4y�NQV��>�<@:�J�i��~e�m�RV��aWԚ<AN�5����d*�𦨩�iEhzݐ��~	���Ɇ�~�t���x����%gؙ>~������ �k�L�� hރ?����7�����/�,\���:&�L���a�3�o�ʗ�L8�j���Κ��-�L���U�Tʻ��D�a����]*�uSn�d��Ԡ��P.鏚,�+Û��N���H��_�*n��S#�������Yd$j�0��cz�I�8��c�Sq�����K�1��Ou�0��l������خ��x�(�>��]����㨏��r�e�:�����Pڹ(#���8g�e��ʃ-��N��^��	����ٹ7vU=��/_�w/�:}=���^܋9�ŋ"xJ��g����������5:[F�Cf5��l�cRXhȌ�H2u���z��:-�l��g���\5���-��+i����wY�N0�_���O=�������a��*)5-���;T�k0�A/�ߜu�N��!��R�,٦L�ï��`�z�S�o[+I�̭����k2��J�	�ʘn �i��۳��j�A�(W�z�qSTx>`�X	�"�	>����{e���O��g���>�A8{�8�,
�d�����f3�bL,n�
�a����?!���$�⍴h.�";���?^�����a#la�i�[<�w22p�:��m��+ie�<��qH
Dn����9e2P��'�,����K-��C� A��rK�j]�o��4D'I9n!���[�n)%���-@(s����D�G�\�����O��`�cʞZ񮯁Ǥ����1��;u��x5�Jz�7T������*`�O��hO�G�����-������GOL���6ޚa9ѿ�Y�I	�k~f6D���%�����#Qf���W�Z����Gx�>�{Q[���/ڎF-�u�ìE;�6��#`��2��(S��!�;���a�,�KR*2?���}u��eӺ�~�r���nL�^�N�٧�V����g�x�Z�����;���Zh@���EMQ�a"7�xH	�p�z��Ӛu/�P�L�0�S�g�ohm��mh�������$�Ű`[�{1|�ՙ"���Ma�!K7��@ ,��hs���) ��"r��s7��"���p��}|�l)r�Pw:�,B��Iv��&�)m9_;5������_�eVTN����!��,
8�G�����u~-�@������Lϱ���9�J�D����Y6:`N���Bt�#Hi�s8�θ>'0�N%]����a��F�	�Wx�k�D�|�9���z��O��"�� |!|���>yf?���U��{�^�g���3�ɻl'�(�+K
tV���c&%���{��E~>1�I���H����� �͇
і�$k��,my���F�5Vڂ44�A���D��6�y�*<u/����sn�� ]k��'�}����ۂ���k���~�ʌDi��lwO\�wdi���ӈ�\� C��L�'����?�5���.�mǣ>ܡ�Pp��o��}��
~�?�}-J��_�5n+�3�*���˳'Ҭy�����NiZSԟQ}�X0
����5�v�5�و���t˧�������p}��N��@��W���2����x�ʱ��~���#����y��g�:��^8��ԍ,o� 	��~b�A��!R�<�DNh�T���M��3�L�f~s"��|l���j�Ĳ©�Z^�5�s8�-��-��pE��Q��R��Ǩ��5*��x�J�y�*�i�u+^��T*c��#��qQ �M��gF��I蚗w�f���ͫ�X���x����Nt�y��n_�T�~����w'b���Y�P��ͣJ��Y��砢�ն�WAtq��md�����T���n<���!�f��n��ۆ4]���0����>���:�T�����!/x8��a�Å�Ç���� #�'HJl5i�R0Œ��2,�8�e�i�I>�K��5	��;Kl�C���A;�֏�v�s�`�h|z��j��]��M�=�Sߒj�N��\h֣��$웒W �-�ƈ���x�m�l��-�t�T�n[�ÜQ4`TO?�q&���N���N_��G����?(��S��V�s`K�eo�ݘY�]�}O]�u�n� �j��Y��]_9�j���	�Nb�.\=Ƿ*��q~��"J8�~܈���37p�0e}��73�mz����m�lR�J��a%Ew*I�-��>q@��B�&H�D�ڦ7�5��U<�M R�+�ѹ��/�m�\Г���]@�V!�z/������l��;�SFd:f��j�k��H���!듂��w���O6��Sh��|�4���C�8=�k�ʕ�j?̯ڋV��/L�~��]D��;����~���B�%fcp�M� V�p9s9�����Q�&@�{�(x0���91a��@��	����ٿ@"S�W�Rm�R���t J�m��7��Ԅ��J���8]�4M�x��|ʽ���G�Fi̋a�,E,��"�� ����il� ���ȅ�� .����:�N�'��.[���y#�#��S�qp>`&߾�nO����/�:
�PZ��Z�$щ!nֆ�p�GěG���IHF��HqV��b����X}�'��P����NA���� h��%����؎�&՝��� �|p{n��lؔ n�,V ��m]�^h9�N
{��Z�<EƪOicR@��`T!���_km�Rn����5�\o��";�&���� ����׾ik���wZ�kX9�LB�w[|,�!��+�7F���ԃ��P �:uv)p!�h��#SJy��,M�/�:k��Kx�n������-*��������6�]�n��j��"���nC�
�F������1�w��@$J��߆��Z6R�KC�s9�����ud��n}0��r>�����]td�U��4xJ{���6���HsVbV�zٰ��z��+ORQ9k��?	w�\UB�U|��ʅ���a���t�7_M�/O���;��$�T���Y��GMFtK:�6��(lW7���sKb����n�Em4|�؃7��h$p��̞��� ��@�ԟiA��V.�B�z�3�����7��#t(+]�J��^�_M�A=@�WneZ2ן������D!�VZ|�!8�����U�w)7'���9�F�W��6A��	�d���� ��$����ܞ��s��������p����y��b����F�H�w-O��_�@~U�C�<�itO��ާD��T���g�'���qL��5��K�ꦤD�툡��M�5�|dK[��@3\�S��7�����q�ڄj���rZ���(Z֞�j��X�u�ߝ:�kհ���h���!�Ѡ{QrV�_��V�$�Ϛ/j�G|
~�ArBg�#	�W�e�h0<��t�$��+W�%����?�������K4f��k�"ނ���d��Q��|7����F�%��} ����ʡ_����J>~8tBf�p����(lH��.�` �6�x�fDuq��H����A;I����A�r�`�&?�Ћݢ����ĵ��� ��Y]���M,F�0 &�s�q���>ǭTx��u��|��y42��\rBs:��'�*Y���+�ތ։����U�>^F�,ዷ��?��ꐪ��ш�!���$��gH�rv��r���dѤ��Ap���d2|�@aJ\t����T�����T~�ٶS�K0,�?���^�C�X�n?��o�@vs��cǥ�ҫZ_Ԇrq~U
a�c4[�&xe���b=�#�5����ʽٖ�*Z��[{]-�m2�Gd��:�D.�\�j�B!��CVS1V#l�F�A����&��^���d�����Mˋ=��pc�Ź�E�<��5#� pM%)D���V.��9B���L�!�]I��)���Z���l��?�s��9����[����� L���gO)S����ֲe%�}��Tf��b+�i]�i��'��E�t�ed��h���k[tE%�6��4��GA�҉�ŐQ�~�d�{�1�����jQ���f^s$k��[��LAMI��zŬ�؀@�u����<����G[��Lc�	�p6
�-���nW�x"u?�p� ��X��1�6_�)�b�Y�Ó	����6�D��>���E��:2��8ٚ�ܦc� ����͙,qd���t�����R�	�z@��M�1è��yzӤ:�|���Z_(��Aͦ����������n;����lP˚�.]���f�a�G�]f=G����Z��d�X�Ż@N�?�z�R���m���rDt�aS���R��'���.��ޝ�7>5��J/�l��ڣ֐d����,�3'�uՓ���{7�T���Q|����B��X0 �q�>�~`SE�{ٹU�x&��6);Em���)�l��u�y�6���+W؎�:�/c�ȹ�eR� ���
�H���PTX_i�UĨ�)b3�`��+*����x�*m׻d�*��X��H�/"����+�;�Wn�r���XF��N�
%�W��K*����?�uZ���h�#+s����#�ܐ lu��iȁ�Z�-�T8�_�9�?�e��;�g�@�`�����EcaN��ң�8����մ�eR�à)�ɱ�2Y����V�O5��`v��)]���r���ZILj��j��Qk���LiԨ��ED������	V:����/~;уo��#YM-
&������_U9+��"?%q����Qd(�M�!�kr�������16T�x3�x����U�~ά�2�:�[F��lr�bH��P�i"��o���./�cQ�^���M�[���mT��������Ɗ�nO�� ���ds�V%ɼ�c�ݿ\�+����s|���z��ݫ2KL��o����r�9o��N���Ī�1��
);���2�a�Qt���Z�cW'`� �����Oo�o�P���DOb|�¿B�Y*���B�Q�F� ���-��bu&;�P;0h�X��%��z���@�q�U���ED�Qo����eS��-�3�{ހf-I�pG�	�	�gG��ئe0�- �f�������*)���	�rjk��z'0h��`:%c�F �m,s
�cR� �"<K/W���n�c�ڻ73��V���W�U0���S���`k�L�G.ԍ-��C �gg<£�u<� =��mE���c�PX��Տ�Xjn�lI��9X�K`�1jἷ���_
�y��p������K�5�p't�R~R	��U�����5�fg���cd��O�g��0��s��}[m+��x��L��7��vb�2C��ku+�����%Y��d>Q�`�y%�Q�~�X�A���a�e���!.ꐾo` �u 
m�)j�;� Z�CQ���,Ϻ��g�CI[���}!P�@`��G�_{Ll8���@�Iʜ���d}�f^$���@���-�D��%����֖���_vl͔�������Sq�;����i���M�v[���-���y�r�-�`��J�l'>��|u�L6>|Sg����Y� Q"�p���u�J�(;޶J�7q�ذSd�����̈́N����&`��Qш��%�h�_�����<��(4/�rrv�sD��k���	��0)���c�%� ?������#��r��o����y���O%�`�>y.��;Q��V�=Ϩxb��aU��^��\�Nl��EA+/��X�'L�A���|���,h��|��#��T�`Gݑ}��.�Rn���Ķ�������
fG�u@� _q��>�k��\��ExȈ���C��
,9~i� K�$#�P
�I�9:����M����U�T޶,_U ڕ+6��>���G�\�ྻ�z��d��mş���l�V�|�G�S�.z�I}!�nu�2k��HЗ*�Yɘp��Q�[w��>�\b;���P�