XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������IMG0yJ���*��M:X���W94ʘ��%w�� 
\xT�F�h��-/r�J3^ם]�Q⩞r���2�sQ@�F܄ˑ����b᪹��^%mҘH��S2����×oX��w�4����2�tIq#��x�^���ʋ�v�2�ȕ?�'ȼ1��,������lW��<�1Ӭn���o��35N�������*�D5w�O�K�57.[�=���v2/��4���/z�3�c�7��	ߒL��͸����!P�9��f����u4u�����M�>��fG��%�))z3C'�2���b��c/�m�G�����=�Wg(����)�`]J���i����绘Y��V�v�P���)?�i��.x�?T5�k�=�6-\@p����jnH�a�X8���C9H��µ��B���ҟW���/���3zb����+o�Y�Pb���������
4Wʹc��\�A{ޠ� u�$]m�n�7H��pK[c����2�/�y'��� ��LR�1��i�o�4� �s�!��S^yPĠU�!`�:�@����G��@T�Oa�� 9���=_<w�vv�����&ܒc��Q�/X�;�������=�6!�BYW��q}�^�t.�FtB��/w�釆.�3�s�.b���f+u����Q����+Q��N� ������O��9��9K_y���#��t�b ����A2�;	��a>(sd[W��Fg�I�Դ��a������K�ηgXlxVHYEB    15bf     890�N�䋙�oL��'Z���n$"/:7�a9�C<3d����p��I����ꑩ�Dqg�\��{-��)ys%�Vo@�x1n��)�����܉��������U}R�Y��p{k��� �\gs��I�8���_@K�l4��0R%ڎ���`o��r�^zBs�G��P)�J�"&ڳ��q�M$)��6Q�Zk�M�~�o?E��JID�CDh��al6�zj��`l�Y���c1kQ��Pb=`�4�g�c���+7�3��ʝiɪ.���t��l�vݰҟa� ����7�����E�܂<c\,����5���V]A����a"�Q�a�m��q h�y��#!W�3�B��A�d��G��J��m��0���'G�Qw�8��n�Y�w�Cg��'ɥ�r�co���!j�ʝbaj�?w������t�O��u��z�0X��{�pp���hGM���[�:`v5tƬXDӧ\��ㅶ�sp6o��( �������*ޫb�V�� �A؆SZ�j���@��2����bd.�*	x�6U8Z����,i�റn���M$��
� �p?�N�T(�š֭�c�	'��ަr�&��>���@����s�D=���6�1sAX^"��Y����z|K�`<_�V��������2�5����[.�)#�Pv�4U+�j2���Ai�Il�Cč�T{D�~rߧ[x�RuY�|I,Dxk�I���$�i�J��63�ї��_�<�K�ǻT"=5��0��m�R��]�×��17�y�^SKV�Ӗ(�} <o�V�s�C�N2`�H�)����Kc����4r�E����������-�b��m	�&�w�^= ���S	Ժ٠�ݻ+*���ZU�
igS2���8�s/��;��B.T7-�����v��:��LK� ���s�)�WR���P{Xx_E&J��4sZFI�KKi������V���^S�AO�S@�]gD)��e$v�crE{���J(C#Z������r���[`��r�+�h;��-����֘�����u�c�u�ӫ7N�hr'�K��)E	%�fʨn�0n�o;N�EP�sE7^~8�d �8q/��z���GY��'��2�	�4.H<�o�2=d�]��y<�k��9`*X��Φ�g�]�q7�帟3�
���R�tc�$29���[�{ g#��J��瓖��&%���7�X>p�f�I�7뾯wLȘ��>�2͘5�
V_O��f�GU6��}�X�����k1C�| L��WB63[&׈�4�P'���($V������p���X~�s�m��N}���$�S� �a7���W�dۘܢ:n�a����:ou�g:4ZCn��)��_�AW�^	��0����g����q���C?��3t���޴�T���f��j���"]��V��xh�̙<c�_�"�ޤ��z3�4J&��DĮ�NuX�%c�I��G�-����t��:zi�<53�5�v%�����3qD#��D.��8ٺn�_��V��`�N���E��`�[xb�΅h�Է�p�s���t�}�tL���#4eA�*�7�b�?�@���^ok��QS3\�n9B��{��-��jm�w�xF0��Q]@*\�|��6�����B��%���k�7��o^�$3ƗĽu4��@���ӺF�K	��ҥ�a�D���2��x���*���_����9�IL Ÿ�)㓝�8Ӆ�KwG#�SY 3�b���5g��V�	-��,�p��t� $���>��׮���p��t*Ѝ����W��X�ST~,N�}o�Ϋj�Tj�?���d�t�CTXE��j�@��Mw�0��y͇_�S<�_C?��2��y���B�{Zj|�W�V�ʝ$�
��^�y*��|��L��V���S�O��§��-m�>�B���k|�&�Z4�h��������Ƣ�H
�VQf�X*��x�NZ��������R$��-]5����	����iޮC�!���o����gN�]x���ad����@��'� H(��6�a8x�a�RlS��ik��G+{`�D��*�����juS��85̐��#���_�DQx&S���㯼x��y+�m@�E���Y�"��ro�]s�r��������S�?�������6�߱�A �b��sW�o�m3u�QD