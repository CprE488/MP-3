XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(�$�����{(�tj��m�u��K��v��Yq��G�6S�Z� �����u�+kH��-�!� �^�Obf0}VH���j߃��`:Gޏg��R�ɪ�S"�JT��[i�P %��eزĽ��9֩v=N?�9^f-��ez��%�w�j#�$ةmC]�7 �J=UHu\��8�M-2���6��ވ]�~����2E�)+��\V����EhZ��:<௩d�Ḡ/
� *#[4:����Z�
���۹�ىu=9!gؚ"=P�DLQO��Q뷉:�
�q: �#��<r/Zq�J�8#�gk�����ξ�OͰ�-O���/H�jXX��\l}�f�,zzo�M/^Ϥ�o?]����M���2?4b����8j�
�ɒnI���D#�?����|�6 2��7^������g� �Y!FEk.����nRb�W]�o��F����Z���ڏf���R(@d���?f�1���|�m��0x�Y-5/T6ZI�P"�~I�u�ٟ�a��$/''�����t)\�&̓g�"�gO�V?�qb3�;$�Ǚ� ��	r2Y�?�<�~u
��4�5�D͋�?fH�Cπ��ۿZ����ssx%թ�5�/�t���Kw'!i��4��V@n��l�"�z 3��`�M�9��\�,ٗ^(��f�vud���΍���0���z� fb�f�3�-؃Ż6��+�C������̣�<X�p��9���TU��U��h#�5N����OArh�C?uL���c�m�}XlxVHYEB    6315    1790�I��-��O2�4��E�R��R�R� �]�؎��p����	y�L�q���&���W=ܴ�ˀ�9h���2�f`����%4�wGy�SD�t��RiHM��]6��Qq�`u�c"2m�i���̒T'I,�#�:��L�������|��%ٷ1�=@d�����t����<�MƷ����8�þ����j);���:~źYX�Ue�f[�#tdAXCȨ@�����1��Y�_�M�.g\I]w��Ǆx��[8������|�Ļ�h�`�!G�n*K�B��t��R�Nk]�6����~_�@�:xJBOЮ!��i{�D��0$�8�*�h�BvŤݎùc�U��`x�-�Ñ�w����&:��@��3�O��3�n�xk+�ϵ�L������jiI ��(񴰍��ɕ�l#OQ�H�1���t�2��t�m�X�k��+�����7�R����m�%��m( o�~*���C��=�V}�N�~gv�o��^�#	fF��R�w��H;��U�Ls�P.�7E�n��W�Zl2��,���O�uK����5��J��0_�9$���������UJ�;�Ik/�����l�5!�|�:*I]y2S	����#]��$ٹ����e��L?�_��jo��m�+�t�ÝBv�Q6��@]M�~�^%��TK����˯���t�`�))���+/º4##:T���6�r�^�pK�ō��vP��Cv8n����L�+$S���ju�L��� ������p��-/`�u���ݶ���In젮l<�&)����?i���812��_:�Q\]:��QT&�J ?TgX���I�գ+����͜`1��5���&��[i+	A�)���>v�����{�%�Ԯ}����D؏�2V"ҏ��8�d�@e8��#�.��΂\���K��qG\eLn�?"�nBǧ��smUa��r#8�>Q��΢'��]�JE�zV�C�[��T>��w0�Jg�TU�ȷz�р
OU,�X�-R�/�g�_��=��g F������o��yQ���0"B�$���a��OBA%7`K@G]���<6��[�Y�q�|0����u	���2o�r�:�֮���ks�H�����"u\�͛@�X dC7%��mgm9R2#�V��7N1�&�rvw�\�����k.��+����*���������ed������,
�	2��M�#��$�Ŗ��}��]�_��ց���o�����SM�͐�~ar��I�״" ��*�{!��ƲTU�]��U� cե'�z �r�(_f|��e�f#�}5X�W�F9>��!�@�l�M�jќg"�����T�H�X2�������:�b=r��I��ih`.%�W�y�,�<�dazg�O}R�V@�*$�ϼ���"���2�T��=���|@��*��ea��^G��REH��6�'M�y��t��1���U���ci��O��i�ڔ����x�:�Z�@�%J���{WG donJ��b������`�EU����V$Y��G�L�e~�-bYi��z�E)���L��L�V#��1��
-TY`����H����[?7�l��.��n"� ���T>o�F�
�c$
&�O����4������?�m9溙f�������G�Q`�6��5��'8��G�-�C/F#�~�l�C�D�,�+���ޗ� `m�1L*6��/���Ax��P�Va,!k�7P7$n=b�8ʞ����_R�=p��t��&���}�C��~�=��u�2*Ї����#��4 t(�JQr�d�d	��l9���5�~a(l��k!K�Ǯ۽���ȹӖ���o]"N�u+E�g�=�pW_�EF0�?+�����h4�,��a�Ռ�d{�4Ki����,
�g�>�G�NgkD��7��/D����Hf�տA=su�C:�,���Y����]�lZ)�V���)Ė��Z����Y��V"ڇ0�%5h�zr���I��Ij�ƚ0���A�����PK`��"�f�����KkՄI��;[�&������{E��U�:�x8y͖URcWsk3�l��eo/������� ��M���\ǚA�=@�=�9|���zəR�����R��A��!]�-I����h�������G)i��̆�Lۀ�B��yh}S�=���u�������܂����������V��[��J�i��ǰ���s$��z�)[;���a�n���)V�0��8.X��M� L|���5B���2����oW9L�^�r�V�)�cИBŕM�R�?�$*b�>s���������Զ2ˌ+�Ņ�n���=��)�f9yx�Ώz�[L_���\qJ��J��S?W
�3.���Kw)�t�V��%������Z�W����ۜ�J*�\EI�4��X�/+M���I&_�ю�W�=[�:{��˃�@��DQ���V�������B�0�� ,�s#;�M�uT��Ӻ�=���� N��Y�*7���*��)J�mM`U-,D��y� >"X^L��a%�	��sFR�fb S�P)C+[֋�%���� ޏ��^.O���Tå�	(�ӷ23�G���OTz$�XC���B��Zz�@4���ܥ�o��gi�:m�2�Z��zJT��%�k[�bI0����N�G�����m�yi��̴�Hn`?Y5�Ǿy�B�V�80��g�Y*�]ӣ���A��V�U(\�^����dpf�W��ÔU�-����c�%������s��BE����7H ��b�K��,U~��"��'�	��fkc��nm�M���js;����v�yD8�|� �QTjkqXX��{{�-��3��]���Zx4
�%���"M�1��h���}��MΜ
��{�,���Lr�tL�E��0�|�&��{d�=k�i�ڗï��+��Т��j�x�w��Z�Z�a��S�h�7��W�8���؂OWq�zH�ҐK��s�%hC��-B�@&'�e�1���6HJe	tb��Z��|�s��jȱ�k���K�0lx6�Z��C> V�8�2�s?�T��Ν��CX�2�ІSl@+�F��O����u�ݶ��m����ւm�n��F@�d��3O��]����j���Iʨ�мz��ZD����x�C����/+.��OW���-�
U���GĻG��3��jC�2����+t��e��mn :�i>�g��w��c����r*iCw`�/�YP�]����������8�;u,�ڎ@>TN��-����Ǫ�B��M	�.��ْc�O�� �_�Ƹa*j����.���{H �<GsZ�@��S/ܤ���x>ɬ�&�EC=}����lbq�n)a���eIj"����|�Ⱥ�d��ý��P���*,_�����z��6��+�'��S�iMN��a>[q�fܦ��Ĥ�. Y��܃�S�F��KI��]��0�����z�8���g�_J���&9^���QCcǢ��1r�^#��[�k�n�s)���a��;1.�w�����<�x��9T�5ݭA��ⴚ-P�\�m4k�ޔ!��9�vz�ĝ�9��ft���D:�+����?X��q9��B賱}��98�R7�1	�����C�J���,�X�F�BOEY�GX���q[�ī�����#y��J;1�2,�ó
��J��'�x�|�������:���"��U�k��]����b�U��R�g��"웟���Cd�M*�m�R�`l��ҧY��h^��U�nV+��,Ͽ<lP�C+?D)$xw���櫗z�4G��:���y�бld�:_Q� n&8��0��%r��^0P�ɶ޷	�{%�����ZduT3'}+y�|�}u�T����i��|������0��[���T���j,Ӽ3/����>�)���EP�.M��G:��R;ֿ�W�����Q�HO췎���@�j��,�)a$p�J���K�}��ezH@���_�r}j_�6 (���;�M4�@(�"��$&�@�s��@�;�#��3\����/�**%Tz��cU1�|��w���y�ق��J
�W��Rtp�:Xv���y�!�j4M6H���x�^���S��q�|��C:mDv�;j�kCUk8򕿦��XOd�M�%*��R�@R]�7(�V�zď���z����������O�Zџ,U$�8d7o���t9[������ʝ�J�n!�k�g�Lh`0�:i��������D���
/e��y��>`�7�4�)�ֿ"�"�bZ��͓�T1�\(�M�>t:$�x��g1[d�Xl�=&�(:���Kd�h�mu&"����T��r�n�0kr� �adkr"lB�ew�P���w`_�r|>��}�k^J�	
���Z��%��*�%~����w�G���ɺn����_��.x�S2�A�摥`�eM|3���-��wdj�Ƀ��"���T:t<'�ڊ� �`v��� ����V�t�^�"^��{S�
2a �l���,"/�S�R�	<+/1UP0ãvވ�m�����������vy{l|.�K�(�.x�Ҿ��Pc�VU�%��:d��A�NzZÖ��C���Z.�p�$kgkə{��C�{���Bx�Y��3� �9�OC߂B����+�\+�fkZ:���#̔����/U�}�`G�����:�9t��{}����Ţ�)Q�m1F����k���!�߼��b,'�X��c1�ol�#D�[�5"xP�~X.�����:�K<���O�_��1jD%V���ǧ�X%cvU�OHwepV��gJ���mŔ��dV�@u�HcH�byù'��߁�a��ϓƛ#�l�-9lH
�$�ߐ��TW��c`^�z���C,�ߚ�\�.X&{ 3�Kw"=�(Ǯ�����Vp���	�����WJ�.�ϯ���_g����O*����n:X���4��r�YjYG��(��o��	�y@�K|D�q��U�DƊ����̊݅� H���U��h+(�q�޼h����r�����2�W[�ba� ^^[x.�۷����ׄ�<~�ÿ��N�Z�A؊ѱ�ݵ�/��ѩ~�x�YVF�(�I���ۆ A��퟿MNs^����N~DV�e�H�� ����vb��rVlp�ZH �^�q��"^���`f�VRL8\2��&ShE2H��s6`o����tQ��g"E�?�����P�k���9aNbu<n�Y��D�j'�Cpq�m��@Cr��&e2��_�v>1��g�:J�q;�`n�tK>+��fSu�ml�����SuSfc�&��B�Hٸ��?_=-w����y��_�1���i[��c^4�m��e�p���ah��'�Iؕ\rV�z��B쪽�{��NE�V����vS��|$V��i2K#n��/�^��c���gD��mQ�]����|L���a���cW�"�B`#˅�Dw��t�� )������誶��0��g�<A��2^�Rw�Vc=�5�I�gui�1h��Q������u�崓���B����~i�S�tˮ�#�ii���N+���^�2+�C�7��K�d)FNjr!���ٶ~�Np��9-*ذg� �p��O�ֆ�MA&1�NQp�L֭�r���(D���GEڜ�̖���^Pi���_qy��A���z�-���n�ݷ4z�?�)�L�偎�Q<���ф��~kq��-��FD�t_�O��=\&�N�o��r8����q �n��hr��!�Ƌ�Zp�{�I�Z(�h֒F6�0}��7B ����������3��R<\"i$sg�����;��O�Q2����j�v�I����z��:�wD�
2��m�f�,��޳��I<����� �W�hq���=�f�t�z������*�����C�Ū/OOU��|��x2�Q`