XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���/��yM�7�Gu3a<P`~�d%����/9̓��3�A���PS�rր����A������~Qv�_�M/l�C�UΔ�]6��"@���;�"�Z�CN�1	��S���h�-(�H!3�	�������g��� ���d �Y��!���7�kB[[���Ĺn��C����d����ʢ�⍝�4OL|��b��
 ^[�Y%e"ϐ�i2i^��o��nѦ���T����&$H�W���n4r�$��6��3|K��7���8b+{��U�Fh�|����^�FS�Lkk��.�����j,�ٷK�A<���@,���3B����{�u�oC�.j�(�a��44�yXcPIg���b��#
H|��r�h̀�?2�e��A08�H`+�Zꂟ-���7Y���55��U�ĥ,#tI��؁8h�lX�D�g�`PuX���<<#�>ʵ��B���,��P,� Ցf�����p0tyuX=��)��~�v_��͏�k��@���B�n��fzK9��=!�z�܍��ͫ1�{�bIyF�frI�:��,��K���ՌW�Q��5����5���U���}�4@�BN�F�H�5���VB��K�f� l�#`�lq�����G��?�ّ��S�H���C!��aGLIQ�+�oK&�6�F����q1�f�e7��'����/u����\�wZ�T�����^�rE��:��5�b�z��[hEJ���$���^�XlxVHYEB    28ae     b60�b	��-~�Cյ���20f� |t�\�ط�Yr�Ot݊���zpE'Y���Of5��ς�:jx�K"l�Bd�x�Őh�}+چ�i�0��9�X� �	I�7}���逝q�k����p�N��!y�}�RG$�L��^<������$|ye8��C�m:'�Hs�9Ep�K3��<�3"1n���3���c/O}IS��Bi=��<����M�uC����O� pf��x�+���U�Yzzȇ �b��X��M'h��f%����.�v�1g�/���3���đ$��r咻(�mt�0��k�Y�� �`���|�j�r�&Ԝ\�.j0� �L�	U�Pt*�4��-a��EI}�Z?1_�\��,�Π#Q
M��DB�"Ygt�JօUD��^LS	��p��h.��1�ޔN����]&��~:Ro�I�b��/�h�w�W�!�b����Lx�*ɦ�KhB��\JY#��c�Jx���������	�X���s{�
�D~=4^�!�\�	�pi-�hL(�"�Y0�����Y"ս�GR������c���N�Ei�	����-�/?q[�M
�\��a��iE�$�B��&$��Q��'tG�f�s&�$�x�ͳ��s��+�kpLz�$;��&�6��1�jU��<���-I_��}:�3�$�8�D����h�Z�����#A�6Ur�Z���.A�u4�	;��w��k�>��vWQƫdE���W�,ʿ���FS
ڭ���5@�s怔�_����i4�x���hJ��w,�>܈Dc���n�m��z���p#�(�:@ˌa����7#�-�.��>��tq�%>󑏯x'Q��4�{��T�>�XA�4=ȟ.�`���<,Q���t��$X"����2��$�ݻv�|Z�C�ɕ��ǣ>-��Ч���p��خZȞam��������_�w���#��	l�c��ee����+�S�Te	�uN"�ω<�=�7�!a�[�C��D#�#u�V-?Jo&2k�AU}҅&�8� ;�j�0�e�4�+�أ7v���1G�*<2�\�[��~����8��赙/h�����g�����L�����[��}��v����p�8L��1�%o�	��r�,NJ!��o����?�(��K:����]17|D9Я��'��/^O�ho"�84	@��F��atUn�&�m4>P��ة�;Z;�[;������Y��d� `�p��V��2�z%�m�bt��.	��o3�.x0�P�x<W^���?F�g\d�^�p��6{wb�)_;d�4b佉z���ߎlVD�No��,��}M�-B깚� �ϯp�"�񐫁ݳ6�+���7D�9.A���+�[*.{�[T�@�u�G2#��
L���<�O��X��?	fd�ؼ}W���+-�.�EW�¸���DOp\�|��C��D6��2n�r��d�iS���_K7=u��nC�r��IMj�$����t��S��~-D8y`Fۏ��PS�X��Hpi�����S���N��㲎��+p{Zŝ�Bi��
A말��^ُ[{Iy�6�EZ��1szް��K[(�ԉ:���KJƉ
�ĿSg9P�9��F�P���:�A��U�b�~�Gׁ�4!��@"�e��FI�m�t��tx���ޣ�rN��9D�="��.�����;��e�4��ԝ�(����w�m�A&S�ď�p\w�E�6�����3a���:&xp+�j�V���ROZ�Ug@E���a�b�5��v��u�}�Jwu�Mw�G���L}�܏v��NQӋ�^Y
/�/����"R�$+&�����X�\�P/�+a�3�L.�Tl�X�D��[j�P����1l���%4p,�55�'�^h��"���\��V��l�d�;3�,`�c�<X�3�Z���}��
y
���y��i��Oor
��Zb��iL��D��������U��
���[�^gv%D�(U��A�����j��M�'T��)�=�L�����~��ڕ�@`b'���^���G��MS��w�E�W3�A�E�p���/��Cq�D�k�������!n{sާ|aeʑ��[�f�fN!i���5��~e�y[&��&�ݱ ���|�5�\��W.�OX)� ��X�W�SSZ���Ϻ�d'�q�w�A8BI���rc^���~��L��������ch��t5Ɏ�eM+�����/,>={5���n�o�~����:0�_���o�i�B;<�3X���~&e�X�Q�[A��6=ˣ��O����\m�E
�n �"%̆����O������s�ݹ��]�H���f���W����;qÃ@Y���vșd_P�M���T�)��>¸���l����m8�}�{:�G���U�е���}N!$��_|q��LU3I��ҷ�]�àu�<�n�T� ������>�Ӵ�X��x�m�8ٓ����2JS��*q�y�缪I>��Vʉ�Xy w����J��qx|#a0�'e��B�ï�]$���Qm\n����x�J� F������F��u��`?<&2����*�&����¤Pa�l���l\����E�@
��>�4��>�������aM��=�_g�`O��:|a!$�8��Sn�)��y�D7K����� J�#�7�bt�/?�����}�z�u��*
$��6��9T"��{��ì$>��s�� �@��H6�?���!��!'�7� ����C�z�����.��R�̕�G�v�ʊ��>�z�xd���+��_*צ�H��cК�/�F��)`8z���D��F��A�=�2ұ�!
LGd���Sd�R}�:/�$�j�*�D�ZiR�9I����:��2c"��k�<�[ޖN�*�p[���&�UN^�ްM� ����+s�