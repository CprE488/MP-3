XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C*6�0��t(��x��`XjZ2M�[?���5����H���'��q�.��28Q���y�xcY���x�H�~;;�xW2�{�N�SjH9�����F���W+ZӸ��R"�J)�51��;zU�˃g�%L��j��/(��D�fߖ!kɽ�$��Z˲�k�i��d�%Rď@ۙ
��gn~K}��!I�����ޣ埼��M������E���@".ǎ��G���N%0<4'K��c�"���Y�I6��]�y&N���r�^rr��ѫh���y�3!w�iw��>j7x��	4�K�쌥48UZ�B��MKz��7�%{/���SGv�_�����>��ǵA9�y��hqܪ1����e�M��N
����4q�/	���=.�B���M;˿QES��6��z�0W豸���8�U)���V�T�0c�eR�k�6 �u�ӯA��fv��k�%��88.�h�����M�}��9�G���\�TQ׈����g�h���T;Da�Rַ�I�-�?t�°��)�St���E�}����s�-0G��ܗ�@2�o6 ��Əm�]=m@[}����K��P�_CXy���(qF�{H�T��
����4u����gm��bG�+t�fTa�x~����g�]�'���[�{9F0+��`��m�������>S�B.������GQ�џ �3e+k�ښF�1^l��&7e\h^�Ab�/5�@>�6�-fdd� ���W|��=4��ƞ�-U����!qXlxVHYEB    6315    1790�����'p"��FlqO*čtb�gn���������l���+���&�3�}�^�cK?=/_�ZH�%s����짘�K�vid+��벳Y�����`q�pV�p*/q��=�x�Ֆr�toI���y˄���9r�3	�Q�0�z�����e�ِ�m���t�/|�;�ј^�.�/�:	��E��4&�	R���|S72�2�(d�����DpmH��=-��'��ЪK��NtJ"��~���pu$�a%S]yR�	���~kţ���o=��+��eJ���f9F� 5!Ӓ����x2�Q���2*zZy
�D�)[��w�|*�6T)\&m�rz�Y%4��@8/VC�"�Ӗ�A��h6,�q��v����^L6��dd#�v�˚�tQK��-��.�В=��Yo�0�cF�02��T$L��x�-��6�3�S5��){��~�B��y��Y/�(���,,���=����Y`�&�bEc>協uL:��x�df��r���x��������x:�<Q�\�"���B!����]�-��%�+���V���tq9���~7'����N������D�b#����ØA<�t\���j�IH��oǋ�{����2�`��o&��?���v�>lS�h%}���W@vk!��Z��ſ{fgHF�R15Jl�3c���c�zvx\\c�!<O��}�0D;������ |�����z#]v��&��Һ U�&�U����C�u��#2
��d�x���r��Dz�_%��o��a�uu�E��Km��g����S�܋W�ag������E/� ����yp�SY����W�˯�IB�4L�HԏF]}9K��ѡh����m���􏪹��wV���O3�2�qI%1,>���5�}����З�z	��O��d!���zOET�w���[�ᖹ�z�'�7yo�gl�|�����r�|��JD����z��T[ .�&d��q0���W�Z�
�����~x��~7�;�g'�Zi+��t��)��T�56f5�<6���V����1��P�y/]BA>��Ⱥ�%f*�d���K�s����R���O�n-_IAn����, �!��<}��Շ'%ӂ4)�P�����G
Y癋�r��C��1mB ��!H�p~�3��-�v��9�n�)�y���� �e�	����A���^.���~O^~ƲQfF���4�qe�~���|���hr'���:��ɟ�5I�+Wrt�8y���|_O�7֕�5ԙ��2�y¾�"�^8m�����m<T��~N"Y"n4�N�y7��P��Nֹ^d� ��50:�JD��m`ж}�C b U{ ��	�(*I�{�_r����kH��/��s'��.��"L��Go��t��k5�@��K�D�D�4Z�+.J�S��ء��'�S�����D&~�������L��	�z
,A>CM8���m�⎙k��Vv[��=л1n�Q`��9���r[���BS�I?۞���f�ݨ,>��)�괔�}��%��l������ ��z*�~G;�*
ۡK_���H�uK��d���	���<L��^(]1�ٽ��S���ap�؃sQ�@N }�8c��b��q���z>������'GA4���A>������Ax��(�?��M��
`X�zR��Hd�r@��|	H�v;?]�:�@I-������S���ً�D}�`��wEG'Z&ۂ?�^��S<���b!�u!ó���+��h���=��K��f�D-��v)-<X���M��y?�� ���x���2���07	 H��VU���\(���"�AO���lc���9�;��C�TF_7���zW�_���s s;_qA��yٱ��&��P�`J���D>_6μ (h��G6����d�0��k��$�s{N����y5:���U,�_�z��>5��唛�	loj�ym%��`;{V��� ������r(�Y���%ݣ�:YRU���ġy����~l�N�_�sz;�Z��Q�k�Д�������]_���q��E񟯶a�����wq��֗]$x�(y��I����3��8��~���%����x���h@������
�h��Qpfc2M>3���TS�3��#�0��o�l�A0����;��]Jh|g,�˂���������k� ���I������Eo$���$��j���Mk���)��EF
%��[ �s�i�r x�@��8�G%/v�Ȫ)�O_=���ıd�."���_�[��7����ץA��=��o
������T\�ۏ��J�u���UگP��]
l�1Q�<�r���.b�7v�9g�r&�3g���V�����h��*S߷�\����DYC�K�y���Ш�8zQB��(�f/�5h{k��Ͼ��N�Ηw����iO��v���A��<D����kH�~�Pã.9��/w7���U>ܞj���)t�,RlSЩY�Ӓxa!#�M%	�fNbmp(/�.~H�ݲ`�)�+b��G��īAa�����V�{�\�60X��Th����h�a:AwS}�8[ɉ	����b����{���A�J��fD�bu��Ӻ��i��cv0�� W<.�n�U�6���'��@�f�V	����d��Y�N[~*�6i`ql���aw<gzjX�s+���< )����b�9�~$��T"a{���$=�"�+�:�A�+��!;�׵)�
M�x���6�3RO��O#�n�$T�0z��d� ʹq�����S��׭��-�=�0�e��Hq�:�7�� A|<�O�n�����5�AJ������+RPV�6�$�I�5S�9�4��'�v�o�y�L�QϑQ	|;|��(�&I}%PX��2w,3�
���[0PVN���M�d�X�s4u��/���L}���}�6�Kp;m��D&օ����'kg2T�0Z�7��}aZ��9qфXw�u���1h_�sd�y"F�M{_�-�%E/��m*�(���*0������ԃ����0񪴯y^��?���%�U#�".�%;���:&	�^ɮ��t�2`���10^$���X8�	>Ʒт�&��!0P�U���vͣ V����[9Bp��(ᐜ˯Ah33�CԲ7��<��_�@�q����Oh �F���$\�]8A\��;��l�`��2~/���s���s�L�q&��r��������/P�$O%D%x��r��}	�ᏹ�z*��Gh"DEPk����e��\��ՙٶ�Y���A�LL&	�K��G�{Q�}�k����)�v�>��n״+��^�$_=v�3&*��M)g��A�}����]J�h�#5H�Q��d�K��f��`��NPa���Ilyj�YQ�v��qa
�I��0o�N��u��i������ڣ>Im���~w0_�*�v�b�9�o�y�Gb���W���{!Z��@�^�ei��o0�����/4s?ND�ak}ﭜ,?O��hm��Zk��Ɗ�3��E����$2�� ��������[�,:i��T��T/ME$�|��n�6����?�g�&/�p:�Mn�^��޳���Fs=	A����uß����Ƭ�)�u�Y�夗<�0}��m*��$)Y�Ν��R�庶E`QCKI��e�!�y|+F;M��k�M�ڸ9�W1/�D�kz��|Ѽp�=���xu<��R�$�ݣ�:%?&g�Y#����fZ�(�8M���>Hs[8?��uPJֽ��~8a�SGq�9E��{��|v7�s�rG�L�n�ZJv'.�bTD���i��l��_�o�)��c���Sd�q�6�/�U��]�����c�h�q��" 4ix^����U�腬J�������UU��ҫ}���l�.�ƥ��1�AD�����!N��k�E�������(���D�讙J��^t�tE���&|~U�9
�b�����,tۗ9Vđ��`�=�B��\�����5�Ô��Io�7����P��ݳ�|�CY{]0(z���ك0��!|�I�R�^-�pD�Ҝ+Z�2m�]��&K�Ɔ�╦���@������Z�Wg�m
�m�m���bruGG�)EdX\4���E@��N�Y�2��ʿv���3�l�8fD����7�jx������mv�a�{���Ԗ����z�f�����^O�;�g&���cd8�>� -��5Wg�2B�t���O�y[�P�4ʷC�� ��rԞr;��)m�eU��]ԁ�;2`?zle
fy([=�g��d+Y�7Z]��)F幦�O	2~�@C�#T�j��4j�w��-�v*�������v��%���{����R3���Ry��-�(Y�`S�˳�&��ҏf�w7��,v�V�ھ���r/�M��!�����E�/�$����pț~�|p����>��
�]u����0%^��t���N��W�f�r�QE�j����e&�}�?RzG+�,�D����j������" Ԁ�������T�K��0{����w�՜8��3���{?���R�q��9��_��� Ap��^���ԉ�M��(s��L�sW�`Fr�r�e�ZzO������F����4��a��wk�+�:ɶ��1dt/jט�a��^���S�UjF��Y#�箏����^������pۚ=�*���.duo�JE���r�=�nO�I��j���A<��E�k��BD)�O��'�1�2�������o��D����"Á.�~>T���Ek�Ft���,�cȃa�h�@�׹��X�D���!�Y-%I����e�` iۅ�"��[SQ�k0(��$~$��p?�
�$�5V��#� `���E�>�������^*#2�Y����L��zD@�%	3#�XQP� ��?�A7��Gt�%�Ţp|����Ƀ��^%���5�K-~2���h�[�n���������벋)D�ta��k�@&�,�),IF�����NAz�D6�BO'�* �/�M��ldT.�p՝�k�g��X�?x�6zz	<��bL����^A�#����K���g�%�z�gN�Xj0��O�*b�c!����X��t�����J�)�������j�`�Y����ƕ!<�Al�ıh?s��l��֔vRƏƒ����j�"�pj��>Tq`V폗	�'g��)�X�|-�,���ͦ�״��"���w��o�n�g)X�	Q�0!K9�T����!��{�Ɣw������o�v��!�ܮ�A�gE���N�R�2�n����Cn/�ܠ�3:\�m�6��B�'g����E�������;�n�
�������G�M��\�+6p����Ґ��>���իB�,�d{�(-��	�Ή޲�����1��ho�XqQ��'�Y�qu���[�Z�����OM��Z�R�5t�r��r&���p����`S�A�2����H��}c]v1��@Aڙ"o�?wt�K���Р�R R���5�U����'ٽ9օg��?Gn]�$���a�E�^�2���Ugo�[3��e3v�7��k:/A������]ǗBt{�����8�#S�y�H|˞�`i�;p��̈���b'�0Y�蒊A�i59�c�-S8����r14f��+�pψb1���%��;��{�ob���D�w9Yֽ�~�醾���NӒ��|QI1����)�90{^�_0ǐ2�w���B�
MpG����dՎ7"�%�/�y|��R�ՠf�M��Ď^}�氦*amn{�XC7�`3.ﾢV����~� vУ��z��<� uS,�Ӡ������i��n����o����Y��	JV@P+C����.L��<�;c{���R��uQ4|��?	�8��b�ll6�3_K��8\�yVC�Ü1�9�ݯ��{Q�r��|!Y��}��J����d��^�#�a�l�NyS��G��h��Ԧ�j%�I9��
!�-�#��r���y$�