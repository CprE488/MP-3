XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����T(�Z��_��{�l՗�Q@�����J6!4�t �=�pr9�?�x���h������bʽ�~i[4��T��.|x�ed�3���}^�?rnM�B���l��9}���LO,���D�/�N*'���:��mN�
G�(�>�� RL�� E6��o9�F ;y�<P:<yܐ�,���w��L���@��j`�P|:(��Nt/j`�Mj���-o���w.{��O�!y��#Jp/eW��`��{��˳/�?�.�)�
ZȍSU���c�:.�M�ǁI��:2�<�����/{��&G�[R~�j�2�O��/��
o�|�V'U=94'q}���C�(���c��W@�oC?G�#�p��8sqi%�ڬ0 v��kO�5����4�)��*�&E�Md��������q�u�i<��� �Qf��9�|)�����{_x.xo��j֜����n�Y��d���˯�]Ѣ����V���<��Aa&�|���?�H��C*���^Z)�=��G�FQ�!���}�u�m�5
�C�іz�V�0/����㮪���]�e��Ms�GRcr����R�"�g{�8<�P�r�C��^�B�B]Kp|f,��mԡ�9yN���dK�0�p8�e�:�����fh��)�݇�w�J�i���X���:���25Ӭqz�!���l�� B�+b���'���>��B'y���>�k]/�H>r���%N�$g�zF,�n8��)/,?1��D��Z(��)}���XlxVHYEB    dd8f    2160�aJ��&V�N����lXMy�������a); �
�\>��΋�3�2AB��,�y$k� N<8lLe���@��Ds�ʸ����T4���^ �zcu��K{\�
��AG���7���ݢE��ì���O���`�Eg����4�y���ֵ�$˾�"��
�F�X�knlߞ�ϸn&�x�ިB���
���m�i�:��$���ٔԚ�E��6$[���v��Fn������<��!=W�ݿ�pw��C����s�D߹����ZS/�_>ݷ�U9��b�cX��F��1�����Gci��=9���q���"��!���0M�g�%Q=�j��Җ��.��ن�7��'q��v�:].6�^Z�J�E��#�ܧ�f?J3޿�ܭ�l�jk����|ڷ��'���:���4��m���5�ڽ�O�gC�F�fU�]�/�QS�`$85�g�?6t�v�y����WI- p����A���2|��B�,�P��h�&�,��H�3-D��R/��V�ϼW`rW�o�4��$�T�
%��
N���*c���it[��@3?�1��t�cn8�4o��ٸ��8�������T>uc���j8MƠ�
��Q�1x�˸K`&�k:x�����yz���ӥ^F����&��<���/�:c���@�$�1o��9'=��n%bC�ʮY�(�������"3�*�'�[#�!��K	Q�A����[o�K��e���5or�n�3�L� �-!���o���K��a�奴�9w��b,x�}oK�P��~F�#0�ϣ�g��I�Lk�(�g'���X�O�A<M"�>2sH��b�g2�PvǗ�G��%���B��Gm��Q5����GG�	є3Ў��|��b0H�l)"s8�����B���n9Oluh��3�����B����\U���>���k�{bĖ�/+$P&�C��e��'����9�ئ�:_>��p�ሷ��D�,ت�bB�BJ����a�t����#�+<��D��u\�
˲�?�Q4 (�8�15�'�M�t�CAu�����sL���E�^>�3�X}̬R)�R�PMEq7�k��s޻Q�\�?��^j����%U�Ub��[w�Z��li�e\�I��N]��<�#��g'�_�(~����/e�,�g3��q��v���}�j�W��n��	@GU����v��_|4�]��u�b�)�~�|e�O�d���@H��߳4�UXV[�il</��;1���D�2!����ĦR�Y��VK����Q�_O�_>U�y�q���m��i��>)s��tl�ƕ.�{4�S���ߥ��V�Z�4�뿰�ӧ*I+�D�it�BA�]��<E�6b�[M�.�̚�@�Y��T�b �s;(5��������E�q�L�`*4���,6��M����	�R�*_�_�k�����r&qeg�Υ�eV4iD������I'q�Q�L�F�k7���׆�LKS`�-��o��?�a��L��x�H�SL�|�y�AU�aݦ%�0zH��
�hB���S;MO/O7�|Ɍ�%�U)[ۆD<?�x!�4A�yP���42�TЊw7ٕMW�8JXi�AT}ʣLu���B]��ZVv���אW�OИ�40L�>��oV��hte<]O�y�?��nȜ$�2t��)���ZWҟ{/�*��j=�(9!K�!K�ȷ��J6{je�	2�c�E��͌��.��-t�J����\�4Y&���)D|��{0�'��8���fH�J_gE���?���jH��^B1P9q�=_
�\w�i頏�1�6��A�r�j����'4]���ƷU����t;p�1h���� F�{2 *�7Fn̅�@�J����z:��#�-,Y�����Pm��T�f�Q�I���4��N�� %��.u������ݛ�Dg�h���,��v�׹��%5V�i�˺3��M�37��9n��8FA��ݜ���Zp4W0G��9]S���W>�Z��~�3*�*IM8-���Z4��֘���C�kyZ��0��֌�³�i��	��q�壶�@�1��엸�Ș����NntJ31�a�-k"�Ē�G��-���5��F���&��X$��&�N�i����_#2�ix���߽�=h��}�G�9�VL/����g˭��C��E߈��B$:g��rd���ƹ�^���ޯ~/�u�ƈ���ߣ��,U#4g��L�(L�_��.y(�x0�#:�����F^�*����u��q�$K���y�z}_��l�\��ϵ�旻o��F��Gɔ�� %�;��6��Tax?(i�W<g�va��z���ͨ��2�r���{��!�гA�"�������ef��6>l>:����_� I(�&`M��j�nFg��x��]Q�`G�8��Vp��!ae]�a����q��ext�kB�/�T��ǜ!\^�6�ѭX�󳷯��{@���t�LS:b'4}���='=���	H'Y�KJ�w���2x��!:��7���Z?��ݫQ��8��"%�Ń���G���14S�KQ�s��(�ſ1�Ҋ LI�{?È���K{ |�`与�y��<?��5��c�Z5�D�]���HL1��W����Z�|�=8��<�ɔy�F����}�`]ͅ+��c�ƒ����k�C�BF�+��D�G$����Q�u��a5N���WHQ�Kvn��m_�z�s��QeG&٤_v�|_=�Ū����dZD���>�=�i5�,�(��]�;���8<��� �%56�S��5#�A)���&�ۀqʰ�"yF���K�U��]���W:z+�� :S+�砉u�˸>Dr=;��Z^���f_ڰ�'"ZJ:�ۡ��-yYNJ��	�`�r��=#���??��ع�C��R�|�M����t3�)S���r4���9]P�3ڿ�v�").����uT��y p�sV썝lq�4��Ǥ�"��10ೝ>�L����N��ClU���hSƓ݃ʻ����Q����ɪ���l�����6,�����J���pAΒ�<�f���X��-'��m�
��h����t�}�+/��վ�.�l�T��E��������S^���!�2�:7���2T�"�i8ś�fߪ��2�Z��:ZP3�Z	��
m��z�播��upv�L��Vf']�`��u��"���ך���y.��A����ͣ��%�F�c��^�O�yB�
�klg��������4��9�1i��qa^�f�U�`��~��bd��&}�qE��9NQ��X��LjLZ��'��d���]o­�+�}P��#��Y����srY&����y���仜/�ޡ�J��x��|��� K�����o�(��~]_dNj���
�/����H�L����A�m��ҝ���T�� B���yřGHQ����8k,�J�A��2�љ�=$�����vc�̷�	@� ��G��C�z	zmR��r|p�������yzK�f�f�gB�|`����^��-cQ���Y���j��^�
���Q�9�+���x2`���%�^e����&�?�mwD�`rL�+��3���<��#����L�����2i�kϨ�a��QmPO	(�e{ڿ���
DUpXY�b���z�E@��Wy}񻼘R�C|��3�l�L��:e	�;[pDH �� �z;�4�Вkm̀�b���(Q�G�~�Ez��'K~�[a#
�.0-ѐ����ԧk0����N7���n[��{�p�$�_x����ڥ
�n

�7/^	��o�Y���[��xU(4ސ�'d�!�����,�`�-��2�em^Ni�(A�`D��O:3��0��'��ͼ#y�g���b�s7>�s�UĠ#�<{��~D/��%>�sL<�D�x�Or,"ҬEǂ�٠��f����S礕'�U��&�O�p��tQ��ղ?�&o l��v���p�������:��c?&Ȇ�I�lL<&h&t|*��:���c|��ng~2�L��NR�+ʌ�ڒ*���2��t�����0�xB;�?�$��T�W�m��A�y��u������E�{�vA�Q,�����יЅ."B4����L����7&Lo���I�)t-T����ъ���%|�ʠm����w�=���u�~�Y� E�I�{��Y����c�w+��.�+��!�sc�~�o��h���0f<oF�\�xڠ(`$-F��%k�|{��g=0t/Z%�S��ǗR�n��	�炑,����8�5��{���<$D�E�	;�Uŧ ��Yw �)y�l��Wz�~[o�hwv��+�To��ǴB	�I�<\Gx����
�ci�Sڔ������b{6o&ӃYt��=[MY*���p?cr���T�+�u�8sv����ofg�b�΃&MƄ˰���εe��R�.U�|5�o��ɜ��x�m�d_�D:Ъ�ͭ}��	̳�	�/1䶺AV��Ȟ���&eX��CM�
��
߶~e�Z�w�o��:a�~��<��]M���eGsP��)��|�U��$E�/����=g�1!L�]︵h����i�(iV�V8l����-��G$�4Uh�L�9���Ht��"�'KF�/�g��K6��l�X�t�q���ĩ�冂}��N��bEO�*�r ��w�U��� i
$���mL�k�cߺ>4[��G�Xɘ�1=v��{����{����b�/۵̰@6�C�����y=>�X�t�ύl�Ou�?�;')NOdÎ�'�$�R^�|ս�iB��~����`b��������(T��oq����k@��V��g��>�؇Ox9_��*ab�.ɼA>����c{�h:�;��j���I�n�2�A����;h�;��bh`�1�JGLxC�|��M����7�Sߨ���Akŭ/�cN4sԦ�'���)�Ðp���,=��ዤOĺ�gUwA�[59��ڗӒglɊLQ��^ͩH�e����)�c}1E��e�	R��Vѧu9D}��ul4>n.��G����b0�����;����<Y>�CR����]/p,@a�	�ֲ}a6�w�1�Sp�Oo��`��e��1�_b���K|ٕp�3y���t�yɼ�T�k�͏t>�w�`n7�*�z����?`e᭼������N���s9�/��m3����'�r^����0�\�0���{�[D�g���0�X�f[+�,r��	�笁Y�����u��Bt��d��c(	g>W!�+�ߔ�e�{T���Pz����E�c��䞖Ѽ��t�8�RP?���N����U�ٽ f��*����z1E��r�b7����V�����v�/z=�q��
5D�x��ps���８3P@����'��C�Rf�;�I'�Hμ���ݏ���W����.�V����贲�6sHk�5��MBM���Q|E��cy�x��^�gC��_-�b�Ѿ���by���=�dc�5�̯%R�{��,�6�we��j[��A L;�I�@��JW��d���Oj�	@:��PLcS5�U��=P7��B&�k, �����(��.����v������s]s*`'�	 �@��_��!6�����w|�Ί���r���7�5~*���E9ۃ$�o�SE�Pń�c�ܰV@D��[��%�m�2G �f�z��i3��Dr��ߣvLz�v��H��r��o�Ă�1���K�&#�� �:���o5� D�!5��#���{�Ĝ�shi�I6ډ����	�u6��In��,�v�'&O�N^�m����(3\�@I��~Y��S����
����äD�n�ZIk�-�H��}Cʻ�A�7�L��LPM�,��o�FV�Ya��Wc��<��ԐE�y�2�޹������;H	IZ�9��/C��k��J�O��\W@@��^����8�O���P�<с�5�c"l���R%X�{��&��c�S��_F��5)o�/���[,V�� ]i��aZ��
�m�} �OI������q��r�g��L��e�%�[�D���iF��~�a�%h�G�6���8��E�n���3�遢����?��9�ʞp!ϹOp%c��3�dUA���,�$��`�֌����q��$^Ae�����vD�FG��(uNLG����yf���"�<l~���1����K����� 5�ޕ�8�ՋD��_�����:��(���7�P��`'�*���?�`Ow�_Hs�X��23
�u��}�բ�Fh�Y�D�����̔go�IB�԰n�T���r���2�c(RD�����rZ�׹@�F�pn����5��:i�b��hVZ)W����U+���"P��5{�Z�ByNY�h6�|*-WqQ�nt��5����đ{����䯤�'��Ec.B&?0Ś��5��k����u93պ��b�4�
i��c�B�?4��r�.�H�/?P�+g��.0g����b�j��e�K���Z��{?��&o��ۡZ4��@L�1�>��4���������.u-E��NL���9sD6N�i�J���P�
3E6V�H���"�Fnʂ!HK�U<6�fk����6Prͦ����9.`0.�W�q�c������>%d[3A�m����`��Ӥ1R�D��	�#�:��9똹�6�23�w���J�'f��8b��{(�[��HѴ�t\���HØG���ݚq ��R f��f@Ox�f� �瓢齁�&֓����U�ㅦ��*���	(��g��59�-��DR3*���C.:�0e�a}��t�{�`�yA
&�l�'i���M��!ﴁH'u0*��/�y`��"�����m
S�<��(�+i�Y^���;:��U��oE5.Ņ�t����vE����r`��y,X/:�-lF���Jm8[U�{�=g�M�,-�|VM�ѠqgZ��ǝݪ���͇��ͧd[���	�۴o��P�;%#H���n)����$�tF$����cD�f)/V�+ӵz�k��K�*0 $;���9sfC��ɟ}])tZ��{�fmҽ�<v�[2�F��>�xRm����M�0�sݪ�N��u��:������:��JpK]��_F=f��-�SW|�:N���	[{�I�����o=wk��#[����k��X��C�iH�r��Xύ`l��<���B��խ���;%�P:���8�w�m��i�
�{�紶n���g|���o�+%�06��(�{KBZU��Cr�āU��~�	ߕ�	WG��.�
����H=I�C�!�$mqW��G�)@^>B\O�v�yS�@FM=,���ʷk�p9B�=���Q�1�_�"�#A׌PK�f�d�Me���r�#�w�4G�äK�HЏN�ާ�Q����`�g�hp��a^����O`���5�`����E�Y����O~R�ٝ1:z���f�&m�7�ig)A���a��%¥�3Y��7����o�`�x����B�T:��/!s�G��|��E:[�W��m	bN�u��?�S�����t��l5�9�١D�u��잻�����V����7-���8?*`��W ���a��Z%��[�������qB��!��ݍ��A u�i�k�����F��*ɂGծc ���P�B���gֈFe�o8$H�pi䙧�<`{�מ�*껗n�s�B�b�`�H��uP&	 ��ebc}2���y���휛e
�0d_$0b'���,G��Ozԫkɉ�]�֊J��!\�aV���A�Z�O��,��g(T<u��I.KJ}�@�c�� D-��|;{$�9v��`�R��D�uc��٘w;ίt)_Z�K����_�
I+��n�����t��`=�v���fr=��4ѶR��	���B��G��ݘ��J���M��<��A�B�bn�@�^�zoNKn;]�G���(o�����'�+��}��9p*l���j��֪��:�B$�G;�ҏ���ی�:A��̖�AS�W$�� /�\�²�����<�3d%����G�d�?ڞ�uٖ��uhZ��y���-$��F�L�������(���M��hgղK�����s|�}����4rƯwR�����᎛�)J��j���ӊ����;&^r֒����/�\(<�҃��d�� �8���d�z���F�=���gSީm�{�z2�앞;���H�Hh�'7����_�Sk�y�����=��Q�]�nݖ��S�vK�����^K*ә!iD���؊�Av��wy��xB/��F���G�
���̔F�z��
ܿ̾����c�$mg�w2�a0�8��:徯��w������"����Lmt�M�
)i����Ż����晸���B��>��O:4�����W�g�0x3)��[�00T �oX*��~
�E܈�@�!�qA��)h���
�����+96��