XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Ӹt,�����{hԇq��Y�M�Ș��w5�|��ޚA����2�����p�L����{�3i<_�Dt2�M=�XX,1^Z7�P������d�IP�i�eX�h	JD��qrmnϔ��Q��������{�=�b�_�Gt�>����<NO���R��lN�p��g6:s�+ñ�����@��ͣ�X�	P(�VD�y�GN��aB�>�H@"���#�X~ծ���vT��f	�+I��<9�4m��"� �=��md�iG��)��]ʯ�&҂�=�O8����-����Q�����U.y�����^�Y�g��,,��� t}'j"���d�O����C�$�;��iK�Ow"���, o!������|6�7�D��v?�M���4�«IY���|]W���`NL[#B���w�c��F4��Cf�T� ��g�/�O�[+lF�[w�gcwg��3#�e.poh\�=�!{F�oS�rl�'�]���8� �3jg�`��=�H[�M�$*�����cH�����*�~�׃u�G&Bt��x�$�(��+�1�8�@v)5	�p=�ᒪ��'ʏ��7���3��𪙵���kb�����!@�������H )�a�/���[�@��2�"����|M��W\�E�`n�\���7�P> w��#����z�uIp�^F�J�����4�M
쵁���5���B�̏������92a_X��!}Z�8`4Ϛ�+�e��*0��f�ke�	Y���0Y��!ҥ�XlxVHYEB    4052    10f0R�m��l� t���R@�����W1x�Su�p�;O�ݳ�R%�5��j�����a�i*U��a3�~��#�Y����M�����G<����9.〾����eD�m�z��ƥ�o[��C�jI�
�vΠ����&��ba���E����(�M�����,qs҂~��
�Wⰵ���Y�=~���8��G?O����Ҫ(���g�D8��a��'{�񵸀O/d����* ��"��(<C O|�R�a�G{.��B�ןz�o"eq�GQ4�K� m����m��0a�ԛ5�(�.�,��y�_Q(U�/9�w�G�
S�������U�p/nIp`��a���w�N�.��n�s+J���Z���+��sXX8�g}d�pT�Δf��`��8�CCeZah�B�u��9뻺Qk�t:=�N ��\gc���|l�Q-���=mt�6�"x�NiX���U�Lʹ�@�����GF	���&K���\ ��G��}d���%��q��m-���qtt�s-�V'@H$�s��������� l@�"��\� �޷��Å���H�m�P{Q��o��K��yI��MD������ͩY]��?�� ��R&���@Ey0֤h�_��m�Y
���av2Wy%[k)����E�m�x�Ee�>���&�+;٬�}5i�m�n}~CF0P�D������KtQ�"Ig�Z����G���M��w<�V�J�6b:P����}����7�_N$xb��JQp��/�	�
�<�""�
[%���A�	0�T�ۧ�^a Zsqv��2����Yx��u:���y%�]������;,fnc�Ęiou}��ad�&�7��cfR�̬iy\��T:��Xz,��I���g*�Ť��LZ�9w��Fd(���?g�푑[�k��!���7�
��s]���w`�DrxJ��!�nka���	܇mƥILA��:����a Yb�<�d~gy3�/G˹�<F�i�E��=��Cb��	&sV(?��,����?��&9aDk-�oLe�(�OmW+;1�`����l�0�E V�.|�y$N�{�����B����g�c����\}K� o+k�#4���%��K�J�����t��)s�/d���%�j�˨��e��?��Wj呰�Xk9y��J#��pV�]�6s��M��ws���������T��|#D� x9�T�i�4ɮ�4� �����b�X8�E�9�N�V{ᘧ��3�����u��KX`�|�{�c)+=�3�c�qO�FN�f��k�ӥGݝq#�=|���Lt��/ź:g�g)>g��s�}�(�_�����xZ�Y��=�)�27g�.������1���f��@����{A��;�x���0�ǆ���ō��SN�uv��ϒ��� �P��a�D$FMZ(�N4
�����'*�q�R�B�Ϸ��2�愘���z�l�&�ԓl�=B8��@Q�����>�:v���=Bu8��Z7w���j�������m%�6�/n<`r�L�7����������5�>xn?��<��`1�525��k	�"N)��.�\>�9��D���ŰV�l��w��� 7��F��¨[�ZQ�.��G-@�r;�H|��t��l
=R����:�N��H���>t�S�N�� |!��h�pFE[�1�'��}�<���s0K����0����|އ%�X/�f�Wm�4�k3���&P(I����*b2�J�y��G��������ʨ/;	��A��[��Vm������F2A���~����-z#�R�9z���+@5�g��As���}f��|򧩹���nr�?�LQH��/Ɩ?����`�?�lm:���v">��L,30�P�e��}���!8 ���*O����֤PX-�+A�����\�������!�>-�5o�P��{��`�1�d,�]%zQ�U��A �J:C�Y���wj_��~�$����/�#����M%��Q�%�lA����Y��������@���@a#c�,}�i�?n�K]�>e+w{a\'�CPD4Б�������-Ǧ>^2��Υ�Ҋ(> ��"	b҉��X��%��[�i�CҢ���G4H<y� �g��<+���:�%�E]U Z��-0KV���T&1��i�U��J�G{�hHb�YǍ�f�@0<8!��[���MPFE��"D��oֆ�ԫ6>��)g�����`}CbY�o��ۥ��_G\4h3%H�X����q���7�y��~��'Y<�[KSU�ҥ�L1�k�P�\*�6 dwNH�֠"?��Q֕}�%D��&��0����=�U�!����Q�s�԰'A��F2|cN2���Q�7z�K�u�ؗ(��/��p�Sj0��Ck��5gcUlt��Ӵ��39��Ъޢd�)T�u���{��tq"���i�����ɅЛ�*�����w���!��j�����	5�E}��d�=�&,mki����2�.M^t�-���*Q���\��e�E��Z������	�A)� `����_�v8r�=h���Д�|b%�
��M{�8a��D����3�E�\|i��Pم���7Nd�����&N8��>�59��	Lp�m�
�X���B2M�d��2c����=E�������vHݯF4`���4��m&�ǌ����l2�1C�ii$ �8K�߀H.�*K���-&|�wf���;�,*M����֖���GGՒs7�9��@%B��`=�
,Sv���ZBJδ��v���j�DD�����PE1$*_����x�9%�bĖ̗�l��������:��UL�\xU�|�ͭ8�%J�JN:k�(>r����u-�@��81PS�t�O���p�~�E��"[5E�=O��Ӊ���G���/#͍p���
9�
/(�iGZt,�l'��ֵ�vD����	@2�&�|��!8�R/e�έ5 ڥ\�R۾�#��|� ����sP�L�|����0��k�K~}x)����m�v�2�;r�
���^����	�q�)�{��cv�sF~��M��n*��\��rP��š�U��/ف��D��%����7�滩��ec[ڒ�^ƨ��L�Gp;Ǧ�RS1��#�F�jf���?l@~��P��G��'�����C>D]'�>��K��y��*���VI���ѡ�!�$�Xx�ϔoA5��eq.�Q�DL �
�((r��
���d�f�NJ7�ICЧ�7K��A0z#EC
f̵Z6��[���,�M�mAer���b=^�L�G@��2F��A�`�A�������|癨�.4�l�dQ[T�8�>UJ�O_Dm��w��1��1)�	ʣ2���?�s�,�NOݣ�J���J���3�<������.&�	�0�7���"���[Nl���);S�;�
�/��M�9�;�2��h���z�Xt��lz�3���L����ln'ݶ�qn�U�$+d�v��Wts���/���5��8���ryO�CL�X��#�e�J��]�s��δ�`�;W�&���SuP�W$@]���Uk-��j�E����Wz����5�I���+3n����?�z�>�y�j��ڧ3r&��	���]?u���N�>�EJ=� �Q#Tw��9��!�]̟z�B��>/��ݨ��ډ,��ڗ���!���0^Mi�6W|���n�{����$:�4���u⪽��%Z�;���uHY��|ty`u{�o����uˈ�D�Aܵ�C��u��J(~o!,�6�d(��y�0���K�=����r5s|N)��*	��4��OEw�Buz	��l���Z�EM�7]�� ��mQx�ޑqN/*�R&w!Kk�'��\U$O
*�Fͱ����\ �}��I�o��� �wt��!�🲏qF��J8���"�p��-äcS�� ���Z���-���i�+���tE�I��+k�m��MUx���M-z>Cu��^\��%E]�Kd	�����!/�[��؁�)�������2�݂0t��̓�p^��i�j���P\�9�����O+ċ�Gt��5�/i�T��g}��A�P���]�:?�@B
t&�k���ʟ�n���
Ύ+e[����${�����1����U-_e)T�̽��+8��;���w��m'	3����2-܌���$�aQ��䳫>熂=MU@�-+5�� �S�?�����uG��;�&�h�2�qr�Ƣ 衂iW�4�J�