XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���٨���Xx�i��'�o�P��3G�mWv�;����ve��+ˋ�#�:J}�� �"���x��ْ��1�~>�U�5���ދ�H��N��I��s�6��+��ݖ���L.���ˁ�t䞆"E�� ����Z�ê��8�!���˜����3�L�gR��$�9�db�l2p���F�V*�LJK�h� y�dBXE�W��bظ�r$��������5���1�;�%�X)I�j�D*�\˸��GƠ�d~�"�CJ
'�U_�& wÏ�v]L��������_M{r>�a�d�vOa#T%Y�T�*x��99Ua�k���aE8�	�S�v�����iH��]�����hFmq�T$��k<�V�d��h׀�r��ӅX(N􊳍�a�~T:����-�ʇ����EWr`�H�¼s]�:9.�b��B�,�@:p�K[�&����ZRWr�fK�eS���J��*�	�:��9�@<�����XxK���}x�,Չ��S�BN�X�F�9:�FS�`.Qa�9QZ�+o�&]r��~��1ҏ��!Cß �w������Ic�B��ߥ������=v�%��k�
9��:nQʈ=�.�9�Ǻ�e_�)�7E�Z��a�ԍ慭=۟���~<FI?G�|qy��Y�A+�t0�h���\R"�\�޿<�'##���)�>�qV>8���M��r������'-ܗ��2���VμzS�B�O4��^���H>�/n�`�����C]�z����ܞXlxVHYEB    15bf     890��"t�t��ڈ��c�ڇ�E�F�;�_d��}S����tP�P� �M�8	Y[�,�d9s|�h��[d��T6���ڵ��X�<D�f`:mz�f�s���FN�?̓GI�9���:9n)��ɩĒ�T>�Uwd1+��������՞�66�L"�1$1[4�n7�n���ƣ�)љ�$9�m�j�
���w&�VU�H��{�/8L�+�� S|�i�3j��:������Y���G��x���C���m��I�]x}gm[�f8MJq� �xOC�����*Q2��ܳ�%/uw�JId�3}�1�'���Ԇo���^^��ӗ(B����RlQ�Ķ�#v(����VS7�NE���W��O"�1��V��e����C����Ek��7����*��4��j�z�ŷ�yv�����AS<�H����>̵��6w@�fPG��G�M��1s
�W��kcVM�{�H6
U�jT;7�e����n}��ݍ����)ߖ�G��`�35�{� Q�;���nx�]�a��߉��
L��ڠ���,@΄v�Z�)S�n)�	�z	�B,يw�[���<:��6�R�'��r��XN���{	�/�
��{�ؑF�ɾ;5����H)˒Lk��@Z������h7]��@m�j�
�u�.>}�qe4�y�H�QF�@�!�S�����ͳ+��s�$]$�ʈ�����wƨ�qʞ�C@���s8%��i"���m�r+�MbY��HFU����N9� �Z��L8lRL,J�$4>9zç��D�,J�$�,�$j���5JAE��;���vgj뵌z2R��;���K[�L�L����FAo�~ԏ[���ȿ!%��'�a����)����77��]�_�St�I޲'����P���J<ڈ��W�IU��\�cw)l�LU��G���/V�E�/r�6���&�o/pq���l
y%�E*�P��^�)�x7�U�j�Q�y��qA.��-�yP7�F+�Ż����%*��Fȧn��]�k��)��	��Ĭ߭e�@ B|�����v�{3�)!����Y�Qt����-�l�)}ȝ�<�3��(׌��"PE�^�egQ�u�D�Գ��3�rx�
cy5��\�XѸ3��O��f�Q�T(0O'�]`�B���G܌��n�9+iA�MW���o�v�޳���*�&>�08��-��$T2L��m6]b�i�O�8-]MP��T�����aIG\".��������Ϥp���dGf��H��c%x�nx���1�B�F�+y&��e�5E�or2���m�mT�'�_�;J��B ��1Z���$
E�d�4��@�Կ�~�
�ɟ2�~����w8���ݎ�Fr����[���Q1�
�n_{e��f6r~�y�h+�Q�{��b_�$��5�m�;�'<��7āK�X�\�j�O#����.��2�<�Q��x��P� �6�X 2���v����pMA�s�fM11�,��u��3��=��0�@+e�j�%en���P���W�0�8�g�ӡ�.Q��CY)�w�ѭ+
�gO�ͧ��1��$͠���\�j�~f��m�W�^K�����!*�"ȳ��5�:b������c�V���3��52��6�ߠE�{ �ۼ�?@������w=�����Ǘ��j��g� �K�l�7?[�M��H�<.YD�f*����8��S9�����Kj2��7��a��Qn��I�Y��xX���/�W���&�V/�������}7}��.� kF/��D��9s� �8>t�d!Ė��:o��iM��Y�?VT�Vo��J@����S_g�E�?�Y���������;�,��lZ4SڪxY/���Y�B�'j2%�g�st��a����͡~�����+�_A�(�He��Kw:���!kMGfIƊ $��y|��֏뉹肔� C��RZ�<�쉬�1�	��rHy�.��?F�:ŏ���f��:O���(�4G}2���"/��n�n^��D�?�{����E��ڟ��$�����������s�f2fexч�b���[=��=��ަV��<�&����1˳儳8y�;h)�E��V�+��
`Y�u�x��#�nEl�G�H���m�R7[u������,l���KB�K����[ v57�: