XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���x!9� ��R�4����پ�ݠT���o�D�]�E��>ne�.��:ܼw�`�E���ޕ����1S�n|\�.�-^�t���������
-@FnK��/R?����c( �FV�5�%�JT������ ���!m1�4�؈B3��I{�.���sI#؍�]}��e�WV��{��9��a/e����W���`���Mr�i��7��snZ��gU���Z?�ʔE/��wL�y������8K�(�"��Y� �K]�2�Q�p�@^P}3����jLk5�MZ�I�<��IMKd8��J�
;N#� p?m2�ߍ����
&+	�7��Ԟ�����t�ޝ�B��;���X�%:ǮN��n�E(�Q�D�7K�ȭ5)�TB������!���}ݷW���ee�~5':�D���	K}�sd�H��AC�S?���n-��2Y�r�^��fE-+$�B��n��6���bjcL��R�+o����}\R�Si}�`�/'�����8���|�nV�r��`�ܿ��-y���ÈԌ���3y^.`�u�!$��~�p�w��IG	�@*)��{���^��t�J�\6��;\!z �!��_��^�6�Q�0��Cb���pL�Z�@����=��N�t�Ǉߗ�~_{��E���k{<�J: S���@�ܮ��-��j�n����3�a2@�i�D]�_E.�}@�Z���>�2��J9����ױ5��]$�"E$��7��(�T�剣 �Y�G�����T�1XlxVHYEB    4284    1110�W�����ț1(��`�O�\�uK�7����e�4��Y�V �"P��)cX)��g`Ʀ~�P����mr0�oO��\�!u���MƆ�u@��jDH�a{�Rԏ'������ֲoR��t}DI�N(���a�n:o�6���W<�ko#�x��?�$��׼T�f��}���b����ѹs�!U����]X粽h����ϛ�1���3�ńؖ��v��%��s��X������m���)<D�j��;4��C�5��>��?	"䊯���IF�ϛA؆M}C���볕@�"B~�8#1�B%ϩ�z��p꽞s�[ �S��Ë�U!�TpŪ���ϕP����7{I��u�h���j�-+��^�2��@�=4*B����M���K>b���hT4��?ަ�<)� �L�y�[��}(�>o�mnNq^�;׬�C��t
��Ws0�m���[�d�qI�"m�t!�=��`���@i�,}��hB�L�.)�>e~�R3q9/Z���%�c�S#�U��(�IAhC�4Ԭ}������)��F���*�֘Q��eK8UA�CĞ�g�.)S�R_p��`�*Yt��>N`
��X����p6K`��,+�w��~�{/:0'|V�+K��\�9�B|0,h����_�2ۈ��x^�ba�=|����9����3=�k�iSu�٪<������-�h�\�y�`�1J��C�я��V�/��Se�����V�o3+�0F����;�k�r�י� �x�����S�}
�,�s���F�!�.���	hG ��N�="�u?OB����{�0���4q��*����5�
	ͿoNG0.t�3HW�b9ϱ��]��"�XN&9�s��l�r�OF{��~'J��������2���D��N	{-`�����; ӌ(��R�����Њӂ
���	���d＇�Z*����<�gAl�T�o�F�)�YP�1AIaU*N9�Y���<�`@���K�lF7쫱�'3�%�y2oYk��4�]EM���H��-R�8hA�-+ej����=y���#��U���|���B�}��y���SQ@-ù�)6���Ǣ$�z�q#���o�ǃ�M�+02Yˤ�U*[Q����O������T�i˩��Od������uM�J�v'��@��֫Kƥ���# pɮ��Q����|3�(�`��5/8%�)����ܗ����v��D�F���^?�W�=-+/�nu�X�C�i�|tA�?�Z���n&���UG'C)����IFH�"�M��I�>�
�f~)�t9{�Z�&�؎|�Կ^�zs)�m�ã�����)�@x�?/�}�z�/T�M�2��h��?�r��w�d�9�GW�V�u�׼����M���7�;7UHj�i��Zet��Rf��`�d�n���Z5�eS��°@�n,��CV~Č��g����Jp�c(�@��(o�|��XV�=8�ۗ��@V�/������y�1����ߑK4x�r�Vt��w�D]�t�}���\r�bQ��X3G3Q��������>����L6�v5�=� m:�AHGM~3����t�Ҭ"~\$��)l@���_?�>�8�-/jGDd6�Ġ4�6U�(�r���5K���l3�n��ٟp N���1�):[�Et�!mND�㥒?tk���鳙�+�����wHzִ�oJ�3>g>�o�(��ח��k���ɾވ�p��l c�I�˾@#ʋK��T�����k�,69e��xr˽��-Wf������6ľ`��������p �� II���;�dT��4�T�֟���}S�p@�u��ݓW\�8��^"n�c�:es!�"��9�>OE�⨮o�5W�v檬�X������[��mk��o�B�&��>}@@��kG����Z��9_WA�����&��J$��R;����.x˲,�w�YOGG��	�&~f���f <�����<�J�@��*L�FS�VC�����T{ȏÕIҸ=��Cw ��X���tF�og�͍���O�|Y���rʌ����E A ݆����ף�#*�O��#F�w��9!'!?��6HH�l+א�2Z�o����g�
������_?��6�Qw4�r�6��t�/*�{Z��9������Y�H:�ҁ�'*���W�-C�Sr0�����M^�:�)$)��Eٵ˴��rB2X���[���C�%AV�ʡ�qx���	����[Kp�/�d�����0&[��u�S�<�d��o�ТD?�<��yW6�s���̽�Nؽ�~Դ6αD�������=(>l������[a�
�>����"����{T�ԝ^iqi?�4�b�V���-��de
E�ُ�q}}rm�S0Ζf����h��舁�JbQ
�n� �^)���,�����hɀ��1yLc.	�[�\����-`@�;��L'��>k%���(��]&1Q�Y�w@���Rʾ��hV��fn/@48��P'	��Q�$�X�Wy~���~�b�l�I��Ȇf�pV\Y��8H���<��Cԝxe�a��,q��xU^˸�	רىyXC{���Gȧ�ݫ�� �C�#$�7��2B_�,(���;��,mن6��O��{���,����U���|.`N"ɒ�(��y��[��%� �~71g*��*K�E��#��s����]�g_�\9�X�,��P��K�h� ������h���ʛ�ELY7�/��h��Z�s���AbIݪ�R�h$~ L/�~�z7��G��%��\*A ���bA5�!,	J��L����~z�b4����~ȶ�Ӆ�9�ǥ����e��U�I�D'��︟R\H9����:���h�A�ѻdE`��N��Sڛ�\	,D ʣX+F^�q�YO��XSұ�L�� 6�����ŢC�J�,�8x��D&���荅��Xu����50-��|y3T:�Fp~�&��f��y�
��{F����ɕj�`����E��+X�Y�0G�� -U��^�8�G��%�)��[��Fa�u_(�p����teL��]�h�k�e��u%��N V��e�+*��9WR�L檪�e�ã��:��K+��ɮw�x���(�e��aG��O�3���9K�w��I���vS����%u��2%����uX�%S�h-hv����N�c��aq�
&����n��3��s5⩴�˱5p��₪7`ȝ��Y ��E}���V�
�"{\��PC	������Mc�;0�y\��b�*)>�D}��ō�)ƪc��79,���`�� t��tU��=�\"e\L�|���L�����ma��0�y�B���Z�ϪЫˊ�^Gk���%��@5JW
{0A�{��[���n�I����F�r\�nz�������܎�@{c+p�1��y���j�I�ЈD��d�]��#�0����V�*�$ K�/
.n$~܋���������G2���ڀ�kL{е$�8�y��{OE�_�	�r���@-��,��A!�7
n!���/U� $������b����4�`g>7�����y}�u�A
$�"�f#�sma�Y�S����o�U�� �W=�{�];� ��-^�Dw�`t�I����0�pO�ހ! H2��[A��E+�rо �r�Zx3��b�ء]��+�C�8��j_��uz[j���STSC�TO'�u�����z�=��B����`�4��HW^TU�����^XR��=n�E^�\�ԉ�>��^V7l�=?Z�җ�ύ���6�6j������T�A�x0�Ql7�X��C�#Ol���>�X��}�j�?޶@�sSL-l�O<�~�2��t�et��V´-�?'��h^�Tz�x�����3�3	w�s��܅��m�O�hm9O[��;�%v�T��C3g���p�H��>֜�$ڵ��f�s;1��BI�}`O���
�����_�^�@�2��8I劋`�8S�.�\I�D�`�X�:-�O��ޢ)b���4��L����H�ޓ���>޿7��̆�9��Ph��o��Biн �-0�,��x)��b�	��yG�՜j�#8m�uQ�?8?GȆ6S�>)�C�Xkk ����n��@��B9fB	�1��D�e��m��>S�2�0��b��W�#��r��:�vMD�����:[%����l%�sp�?{��Ԯ:H��)�X�þk�`(xPuB�8�k�q͒���רFu�3%��9��JzwR%߲ދĮ��L�D\77¡Bf�[�����fʧX(����v