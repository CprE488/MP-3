XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����y2U,�8�:�1ie�m��9��,�}��Vcg2�N��n�H�|	�}?%nȮ�Xi!��Z�)}�-��KZ�C`��R��*$�z�Z���o6��&�C��@�]a�*<۰bj�g�5���H��EF!�g�+��ye��.���A��r+LO���/�PX2�4����19�*�P5�&��!]�A�; �n�#\�l�\�]_�ė7I���%�O��Bk ��C�~k�Hj�:�	!�Sb�4Vr6)���f�*������,���� �������wJ�/�ث�<t�
�����(ÒI&�BxrOž �31:Dl��2U��S�����֍*_"���&N��
�}xj��O�6"B���ǀ�Ҷ��,�_[����ç�����`����0 �h�����ޟ,b�� �C���Y��,�/C��FQ��}�����V��:@8$*���*��� �=���zzE~:X-�y�f�S6cx;O����h4��+��iK�}�L뵬j��J%6&2���c]��Ɩf�;x�k)e��	���?�(1{���������'M�n��&q�݃��w��t3����@Z)�.(�-!Dk�$���J*ж����`�ޖlV�Q0D�|�IJMHJ���ZжG��hM[BM���i�q��BT]H�n�\x�jιs���~��֒� �hʳ�`����p���`I9�A�6��1��7�R=�n�(rL82�{�����/V%�	������XlxVHYEB    1a34     990k�t�76C ��{�	
�0T*��r��h*d;�k8�4��{K�p0�k���	'����#s�bsj�\�;R�LYT�-)�j�f��TK��E�`z580�z>x��k �ȇi#����e������_�'		,T�o�*���t�Nz'	�z�.0b�G��6G��J�u���W\;�OI����5� 5�����K��u�5�+��n�P�����c8.:^��k�]��J�v���w/q�qਥ�K��<�{�RG�w�k��2����.+�Z��V��Y�f��p�6.oU��DG��#6lh�W4fIU��е��0�9�մOI�&k`J�Nh�\s��y��V��PP=����B�#n��]�������R��T�-Z"�	��Z�Zٛi�f���&�Ӵɏt�u��^�Ԫy'��3P�
����v̓�"��c��32�$X�쓜+f�޽r�V��D��
�ns"qb�0�Ɍ���?4-�Q9���\u<!���g�wz����B�@ w�*/M��9�9�s�C?�/}�*y�)���p�����c�4I��vGS֤��t�x�  �#m�T�[�˟[���D2O�͕�\<'��8/>����<,~�Wc!�4vh�W�]n�� ���,N-�"NC�>oǷT1�(:U�����F"�j ���gu���
�͎�8���W�HW�G:��dӲn=�;Y"�<���RK>s����]P�*V�Tn��Sy�~�<�|����h�gá�(�]����e�wϊ���\�u���#�E��������5����L�mm��� �r�%\LY@��������5���b��̍���~$����BdXk�Mig�%�LV>��[a�v&2�W�%N��Db9g�縀���40��^�h��#���Sb�_�������"E�}8��{�<��=���vl�c	��9��G��ml��ͨ����b(j��V��o?���a�����]����@�7�����B0�춳m��1Y�X��D���<8�?�Bʬ�N Fa�L>Ù"�j�6���kw ���,�k�}Bf���q&�5ʺ8��F.��}�r�!8�&2US	`9'b�,�����-e��J;fB1�N���YN$QgFoP��~���w��
?բ���`$�-����+�"�B�"�<S�Z5ܟ�a�H����"`����{Tc�?��Z���3�S\B��"�����,P��..���䚧����Ȉ@�"DZ�`ב���/So��������y��7��o8�P?�.%~]�"{������e������+�έ���,��9���H�(�{��+���)}\֡m��QԟPP��A<���|I �+����:�w^޺\���d�_@��J˝l�Y��t���D�j�iP��Et���8^�%��7"�g�Ţ�ͅ�]�/)W:./�#k�G1��U�׷��OXa9�c�]��������gzIʭk�ȇ,��"�
2�d*.i/���ۈz���T�g0��?��vV�6� �'	�>9�\��eRyj2�l`���p��Q�lOaI+J�/���Uk}Y��>u@d,���6�W� èk>!)��	� ؤ���˹"RL�h'1�N�3�I96b�&ڰ��xF)�� n����J���6�RQ݇�hxu��Ip��%�'V2��9M"z��Vc�y�:�;��gٸ-�,�U��Q^�\4�+��O^�p8Oᘘ	$�ST��E�N�r+��}[��q�[�'��w��x�d�ݿ\3F�3�i����'�P�v�6Q���0���UY}$ʔ-��I$�[UҶ��U�l$xh��37�|��,������?D��� �:�k���+MK��x���i�����Q�a�ץx=��4>�Zh�S+�(tUy]8�6qC_��$F橝���;�t�^4С�/x��S�����H��M�lTR���8�g��︘���l5��-P|L���������ds��7��tbŽ����T�Mpo���f1妡:�e�QQ�)����~��vg�����!g���R���]pѺiR�=
~�b�E"�ڳ1�]����EB�<��R<�Jj��Ei:�1׷���$����ܗ��Sm]C���G��{!�G1�"�^Op�Y�Xx��-/Pb�i�������\��UC�!`)z�0H�ic24�Ԉ��qO�����v��7�{�<HԻ���-P��4�Z)�d�pY�kM����OiC;OsA�*n�d�њ+	�������EyJ����V|�����F�WS܈7�+P�D;/�lZ�]����~��<�Vs{���,\�V��3�xn���P:�wn0��'QVcs���+�ɡ����_<7}���DG���K�Ȟ{�+�Y�B��~W�$�g޴K���w?i(�r�