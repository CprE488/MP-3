XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ډY� cd谏��[�ŋ�!Q�I
������ {�_������ �"���q���AQ&sɲ<u��'@-P]�a4C�\L��Q^>o`���CV��j�7;�B�ڂA��g5��Ve�%�ĩTc_%�%���¥��J�҂(�+@�F:W��>��~������#��y�[�a��TF7�~��_{WǾ�6&
B�㠷�e-�S/-(9�:�>D��*��eDg{�Rܹ�lr�+��22�-�w">-��k]F�����a�X��u.Q*���,�,pӞ[�9�FZ�c�x���]�x{���x��b[��k0
tp�dO>�&y�����w�	�MѸ	];G��{s�g�9TI�Y�_�lb0�\��)@�v���Za�b���MF�a��;�� ���zlY�H��Ӕ���s����F�+F|�b)��.�=�R�N��0!�GW�ƿL�p��~��"�5�L��A!�m$�zx�����7;jd�Pcb]��$-�:<ryxG��Sek��e��Z���(ܘӆ
M�j;O\m��z]{�kϯ��k-�D�t=&�eǧ/7�g�L�1N杶�U��L�"�2���9��	`���*<sl`�������l��v�qc��E�A-I�
+�V��s�rا�n����a��g�Q�S{n��S*�҃�kd�Ԝ$0"lFvy������O$ˀ3\�~�QEr��.���PTü�T��~Sg�`u�o2S�c	�G�nB��T�%)G����Q5_��)���A�ǝ���XlxVHYEB    1847     900ݬ���a�k�2,oᑊοS����)�@|�а[��>0����b�/�ρ'� 8��\���W��wi(|���!�ȿD	?��@�q3��Lae��_VW�R'u;$��2�bցd*X��<�98�כ���Uuϵ�{C�v3�h�vd���𢡄Sܞ�p�Tح�uJs�PR�wma��'k�����l5�4���"}K�����u�P���5��Z�\KY8b.z���T��TH^i�麥
hbo�D#��B,ąNI@�m�hQ+�ꃦ�:�9�����&�_;��f"���]�d�~ԡ��zl@c_�-y��q����5�@���]��,EYZtR�s4퇎��$�%fG��N{�!(�9��߭}!!L1X���(��g�nW�E4��G��:�N��y��]�	%%jE��׭wI�cCVMR���1�>�ѐ�jo'ZtU�[��f���OJ�D��\�'ƙ�;˩�@!i%�N���i���-��W�W��ʎ'��o!k4�����:��Y%�#"���z� S ���	ZO4n5�Ȩ>Y�M�x�P�'e�M!�t�����H#���u/��W�����'���q:�1��	wxVq�f� �֥�m�azf�Dp�4��yuu10��P��B'��l�:�����{�ǘ���;�,�vx)5yű;�b է�0�T¥����
����Y�G�[�Q�&u(]�T{��!���D��*���)�R�`v:�۲�m~m�E��N%���,���t�����6j��͊w���h�?":O�_zW�2�rr��±���֌Tq	�����j��:a��7f���d�WgwQ����`ke������m�?~�L�b*v��3�<�~&X{�c$��n�T{�r� �Ю$�@F#�J:��6�2W�0[%U�4b��׫SC1�ٮC������gb��� ��'7�V�*��>m��g�$�a����#?Ѽ�)"����#���_�,|%h��f�X�lu��fdm�"l��4��F�/9�DzO5N�< �8�����\�JĞSc�Å�))�z���
���0�4��$�<�:f��H78�ڞ>0�MU����%Ǻ��L8��q�r�#]��[��ُ���(mhZj�r��s�G�]�}�k�%q@+�ˏ��n�fC��y`j�ԑI�+?E/xR�L��b P�J�؉�y0:�����	����Դ���L��Æ�\*/�Ao�����+#�3���)<B��o��}�<���X�_�ݢqt� nZ"pd3�jb�娻yi�����3�������L��OC+�_� (
�"E�K9hd����"C�Q���Ձ'`��L���7�ԷRgq�?�+�������g�Fr��ub�c=l�TX'3�aя�3�M`(X�nܾ)���#4�.{�Չ$L\+�nG�4�N˸���?a�%��c�
6�����_?���=�*��xRe�K����q����d�Γ�Q��Fl���@t��*�a��*�����Qv���$/m,����(;�eN����4��U��MB��6���iݕ�5ߧ4w�֖�m�12t�Ll0��W�&)�W�-$iH�.�#�lqt�WDVn�����yi��0w�u�@Rv���s�Vv#E��I��kp�<�^������ј '�m�O/��0Y��OAp<�7;�N���p�/�8�=jI�L4`w���[%,�t���Jm8&�Be��5�1���<��Ť�ۑ�����}�"���w��GH�RXR�4���1i�Y���
�US��>a�%�{�����`�f���*0v�x��� ��7���TR�=�-Q�˟z�����ǹ�ͬ��dn�_�0��L�ўOOT%�������� ���1�&�_� ��a�3lhK��F�9���>�g��L�Ь��c�܏X�{w����������&���¯�G{��9��cU�b���,迦��#`b�P���������G� Ī�[\{������Ƙ2�q�e�Ę��@&���i���Svr�n@���Ά%ʦ&����b�3K��7ԍƈ)%>�x��{��m�^5�{:.B�В��*�g	|�C`��]�(�P�Q-��a�;��T�.��RGkh/^�ȁ�+<ѧ]�-�׻ �S��ɖ���^ÜPjOj>���ӽ<	��A*��'�����D�$)���}D48k�ض�'����az)Z�T���X�ZQ�2��.�j����@�[�$ʏn�^u�Cʱ+�ˤ 4�&�X��Pd��{�/���b�l�c�"�