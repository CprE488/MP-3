XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����6�2uҘ;y%D0��������L��?p�;"^�-k�d�FXǲ]�Y��=�#e���[Z}���TE�YMF����/e��P�Թ�Oլn�r�m4#(R A׋�n�'p1��[�}<@m�� -�<uMD�p+eK���� �ҫw9��6e�r��%V��T|k������Q�a��F��bC6�?�&CE��suw2� ���ɽ�_|մ3!���#�ʱ�끪T=M��k	�`�u7�
F@���$�O�c\�I�#�DAL$�S]�q�Fѐ]?a��K�4�]�䪈={�+�&�.8�rb���V���Vi���㉫}]�˙.3H�eNu�����f5Q>�LT�I�3���
�O�*����ԍ�Z��kM䧽���U���,?�i���6�[3�������#瓄N���/w��n�p�m��gKJޗ�@�w#T.�p��.����G3b��}��`;�y�UaB{ޝ.%�F�s�9����R�k��D���2�t0y�4z���uFx!�:ue�C�aI��0�9�p���o9���
B����]ǯHM7�H����vҿ����h�G�&�
�F����&��i	m4�Es�_Z�����.j�A��[�G�w"�������̭��*���Q-q5;��9
w���XYa\`�~܈�B$5:��E�~�;Ǎ�� MZz�;���æ4�ܢh�X\��M������UZs�06#	Q�;Rٓ�t��eԄ2�)�<�5��2�J6hD-XlxVHYEB    28ae     b60�YX�(j�i/���E��9v"zu FI�*Y9���5W��Y��͠=�A2�Rԕ5D��;��T���EKM�//�Fw�0\�%\"7��5:j��gx��� ��j�����wf��8�F§�,0U�͇�6D���bx�O�cG����2,l���&OC���",@$3	������v��&�sOF�͞�@�В,��o�U��u��.�9����L=��*�Km��͈()	>���{�Y��	����p����J�b�Y22>��`;pY�ث��Q�ݧf��aE&\���3���%ɔ6�4<`��3R���{�3�b�?uā$�iF@��^M�J�#EOy\���@�Fe���U&p��>禡���j�3�<D_ЕJF�8C�ofm:*s�J��?��׵�aA�W{M�O��6^	E[2�ځ�J�\q:x��b�j��a+�B^W�Z���
S?�� �ي3�R{ɋ�+x������#?R6*.���	���y���ȍ�W �E���7Kz� c�E�Pȫ��F�[��F.�*�!"�%�M���octV ���T�ȿuQ���
�,�J�g`�ɋH63c$����{b�ȳ���¥\��rԠ�h��<�3���-E�e�|�rv���IDڌL�I=��#�NFvD�"	�4���N[�V���Q�n�ՓGXC@48�N�E��H�� T1/lI���2��E���PSM���Q�5]�@�-�WaWO�эJ����I�1���O`��� � ��	�v�9�`/Qw������#�bE��9�F�"��A�S����ц�0�:�r�R)�5~:��Hx���H�?.+s5톾dlh����-�J�CK=������{�Hf� cX�c�7j�ǅei5*u��v:��eޔרw����|n�����0Hc d�u��!�pJo����N����HMv��+s�w��v�۴����U�s���ZŤ;2�����,S���6iG������>�R鵕��1�ie#Y�j۷qSꚶ�dm_T���?Ӯk{�]
��èB�А�Y��yW�3hrxE4�c1�N)4綾��^�<���eӽ=z�b���+�փ�t^Tc#��ǖk�YU<�bj�����>ғ��?��&�A�x�غ���m���K|g[t��>ȟc�6�����s�t?�8+F�ey��"�� ��sty�p������uD��0� ��-��y2�M�]Y[H�nk�ѱ�6�^�Mی��'n�����ܨP0�_J��}$��ƾ��͸r����� a�������a�c�@j#��Dx��"�TF��^�����XM�,c��.����;`:�~q �rf1��ޓd���tB�}�y
m>X�˟6�g��X�����ͳ�Bmj��F�ܩv�g6W.�l
�1��Β�Lr�Z0z�^|�*�K��E;1�ҽo|�$El�F
�\[#ƖI˫Ɠ�p&��(+=�������,t�_^%p�F����o�=� ��p�⻯O��E��5��4�13$H^9���a�D��j
�����������QG��{���j�#z��m�U-`B�"��l��ذ>OI騜���"Q����f�/\��p.k|)J�=�}}&k\0X��1�0q���%3����HVn{��M>������r��'�4����=[�I��`�fF�]�795�p��L��2�f�`� �S�݃���r	-�;�x�T/L��68����	B�\��:���pzϡn��s�gʫ�:v�h���oU�%̝[w�X\��W ��� I�Z7ql�p!9{��lDn���8����;s^9_����P����`�N\8��ʨ�Y�𭺺�����nIu�~)�����j7k7���"b3��;��Q���t��-��-�uՍ%��Ӕ��g�G��DZ>n���GC9_B����g�;S����C{����6^�+6ݻ���5{�>�^��V ����<��h�	"��6��HI3����a��'�|%V�N���o��`p��@����zE��`cN3��0��7�L��^Cz(����8=�:��$��f9�ƗAvF�w�I��:r�������`�sh��M��+�j��^��*�u�z^��2�/ck�$U�orN�Վ�ͦ�L�-�,IW@�t�%;c�NOZ���{\3jhX����nܩ���L�k#b�o	���J�;*W�MH���}�����+�L���p�ҧ0	������1���B�&���%k�A�cş��!x�Ӕ���z��<��UB�>A�D�0XP=797VpZ:�G���]l-��`QoDL�U�k��tr*4�+��r8�R� �4A�G1J�PW5S����OQ�ϡ9� ��L4k]u�)-�0�	@!����X�2ڥ�4x�a-�>�nT�,�mq4�x�j[�p�q��W޿Q�gDbq��K����(��z�_g�՝	PCK����3��ͯ^Se#s�7>\��˻}�����׬@��P�[�4�i���,_z�//=��k�����I^7��b�]yV;*4u���\������M�����|������T���E��w	��
�ET��u�3��0�'�u�� (9(�%i"L��?���ek'��#3����� �Ia��Z�;g�j�S���Xoe=�=� �"�m�f�mA��S�TZ���AF����i���q0����b[��:6>-����XI�!���V�qlA����/�ī���ئ>g�<}��Oj���4��(����l��*��ۊ�K�(E���n���awWX��>��v��g�	��S����ʆ�w�*Rw1��J�A���]�B2�_��3~�