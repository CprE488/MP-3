XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������&7D~�I�?�!m�\L�����U��Ys�	�]�c�TXtN������?N̝����g�2����C��<�($��1��Cj��	=�U�� Z��Rjx�*�FA�k���f}c�ͧ���n�K�.�(q�{��ȗ4�ZK �?H@��	����i�����执
��}���s�k>=��c��m�ǂm�n��]�[jr�〾��������Kt�I�!:��^ �vY�9!�s�&���$����mԶ�|�2��]8����FVK��ݹ�`��9�HW\m���t9'ưB�`�w{-r�[Zϡ*@��L=ŵ(N<%T�Ś!p��c;�Ȭ��$�'nΰHAՇqC%.���LQ�IDJ�f�����	%*;�7����}Ϭj&�3�'4��]TƧ�[�Ű9���.�ʃ��t0[���C=b�s�X~fe���s�x{�䳲�-`���N(�y�#3�/���6������@Z��Wf&�����y���)Ë�wYzNk�|.������,.u`���'��$�ƶc�Nc}m�=

2����8��Qz�g46�h�Ɓ& ��RW�8��}K��bb/�����-�W��0Z��K R7��^w��P�X�Z(�2�%��	G2H�[ݧO���C���g2�K��>�����e�*�`0��wv;f��QDΗ�o�5�}�V��Mޱ 4x�
ʞ�?�y�3Y�,����3�O��x-��x���(M+�GXlxVHYEB     f9d     6c00c�����$�b��zo$����| 4�J���~��,��6WW����A��zy�����p���R��ka�iP�E�!���fi9N�ߣ&�Y$���?��/�R���N�^}�,K�k{�^�1�NLMܒ��:�/"P��9�w��.:(�IZ���ƫ=xH~��*K
 4��j�B��(��ں��i�,<쫷� �n� �@��/�Y�P�����Y�c�ʳ��aR��m&�LU�R��C�����c�Ub����Tb�E�pd��m}ذc�r�/{����'�b@K��ْ�Y��Y7���ER�)u�XM�^�kw��5)����1:~$1���0#����>�<tnո�ЂשA��H��\�ca3QQq��Vu֫n@��� ��P#��~9+9�;S�ar������`��v+�	z�3#tܣ�%FE�l�0Px���s�O�tBk�Ȣ���*����A`��Ƒ}��(�7��_N0���@���,�����>)ȿ��L�%��D�/�aB�S�:�P�[��%�]�{��M��wc�tc�Q�e�����H��C�Y���1�ν��~&�q:����l�`��eS[la�1�'!P1`���s�S��H���Ŭ9���/�9��2jQL�N�I�eU2�d�������z���(���%���-��O�7�z�����)���I:�I��$��ٶ�E`6j[�˜^���}� Y=�%nrளjlfx��-'Y��粨���u׊�,����+ּ�l/�=�ѵ������FWT�ݮUF^�F���,3�H���bW���3ȹ.&��ts�
���r?�F���ɠ�Y����g@��G�4�L%������ղߎώ�YN�yB�S��}��<�>:|5�u�'a5��7��.�柮
�}r��Jv��$|J@Ƅ����/�r�(H���98S�����iO�W��X:Pr�����K~�*����HB��h�߅{�����v�CR�����YD>S�ijf����E2|�d_�--!뀼tł@'�gJtN=Ȗ5�-]G2�G�~�}ϫ����ie3S��;��a~�|�Ғ�����}�mE�	؄���rs����fԯ�uQ�@>��5���U94��J��4�.�I���y[+H�+�����j\�Ϣp����kh��j�k*�Yޕڐ�|�$d�?ۢ�6ҡ�򏉌�g�7x�Վˌ@�֎�����k���ؑN:!CS��М�Nu�6����jJQp����l�z:521y)Qq��OKN�O�⎲K�<��b[z�dN�@���M�, n����$6a�k�'�_U~�TkR�}Fk0s,z�mC�C������[v-�'�sO���i�bZ���[P�a�Ws���֌>��)+G��y�O~Ot��o:r��;*�)�R�ekq��iKl����E�adc�b����4	��@bw
�:y���=NU0�^�B���Mt#v�h͜_�� �����e���~<����O��!� '��D��0��)�k"�[0�]��彍톷��][�si�DZ��˸�\��50T���J���\���%��QT
�n�
��F\�iU@C�u����:�O<,h�C���[{�x���������Z�����l��� �TeQiei)�S�β)�5Q�tïtK}he �r'��]��������j�'��]�+�k�G���F��yWf��c}b|�c