XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&�x�x�wl�qAӾm����=tQ��-P.�\���!�0�WB����y[�a[`߂!�\o]�$�֞����7�C{�B�MMW�Vu�h���׫�|�Ql�	�#}]��_������B�D��7�FX2�SN���ya����Ħ������B��N�Z����4j8�/�T;�|��:i��a^�/%��U�Y�C���-�q������z~����tb:2��H�;�H�ze\�����f�`�V� r�"��a�����Lx�N��^�\��^�KW�;QR��Cb}�?�����Oz�a�sl����v
 �ٹa����v��x�b�R=y`�אR���=�ߕ��r�)P�g�i��L�6`f	�UCz
~�MVhA��`�Z��DpQ�xtby@U[d= x����w���iϗ=���դ��)�1��iE`��R���`��ڹ0�b��/֨քD]G��֬��,q�'9΅�BT���6�>q�h��&��Ԡ�&n�a���~2��.�P�C�i�PD/S�V�G9 �ʉI���w&�:n,M�w�|�Z]�I@(u�t���	�2`�R�Ms�r ����Ek\l���M�Im��?�28�#نC�\�L���I��:!U_~E��I��ݱ�K��\!���T�Qq�nƒW:[7�Ex�m��eR�죸u9�R���/��UC�gF!�C���[�
z�P#gw�p��ɚ��{K��=�*^�[>��[�,���S�T�m��qC�YB��h� *t�ކ�!XlxVHYEB    1448     800C�j�$������6�Y�,���
�M���u+J�/�)��
�X{w�+6�Y�uP x{(.�x3����j(_�2���F�o_��T1��;�	T�PV/[��Չ���W�ݯ̇��X�Q
��9B���ֳ5T&�X��5�A������8Ն|Ou�2)�*��*�]�����Tc(�.�W(rq0��|�*��8�� X�^��J�+Z��!h����w�	d`���������5O�_�p�n`[F-T����#�oY��Zk���q�UE��0~O�~*���?�9q5��4�I_�1(�:+�Uؿ��!�����;�y��\��d�i�z���(���P�58,I1��n?���i�Ts����1��?L7�]$=#AdBǝOQ٢<�ջC�ބ�Tц�Qej��ܑ���g&��w���V
In�B(� +)�� �\��͇)+Xt1<2�MIf�c�v62��qF��=�����Ц��[zt@�l�d�=F+Д���M� �t �q�<���um�=�A�e�%�h�f&����j!ܸUE�v2�%BlP�.�9/Z���N�e�����bq.�\2ѭb���V�S��������d���M]v�)��V�v�q��n��4���7��z ���r��o�N��L��}�@y��������Z�B���_�4iAh��@��$ݠ��(xd��Ŀ�s�OJR��ʬ�Ɔ*�*�l"|�jn@�)�jk�����3�I�;ۋ������ρt�)���"�ݿ��X�������ã�ɺⴖ�t�j�^J�LG�p��v,���M�Ƚ�M�� &g��#�L�Jq%�IÖ)]��`���m�<�����*-����f2F�VeO���s�2)T\�����0x�f�wt��c�tu{e@z�z��-��c�f)$�U*�I�i�ZB/?�����d.<B�:5����@P�
a&���׼����J��	���:b�I�iv h��N�Q5�����&��R�K#��E�&�oФ���mG�������֞��S�E���>B��]ķS�'���2Sdp�;�.Y�_��v��Ȑ��e��;�I^B�;:N'�WQ܏u�ǋŵ���������䆛2���V��Ť6E��2��M��V[�g��k���Iu��/^�O����=�K�$0QK8qw�R]d�����yT>V�8Ç��ԗ]��.�e����	�q�έ$�D�.��?[�O�nT�|���� �SB*�)7�ox��w1,�N���n����t,���s�.-��G��N|�2d��&4��l2	-Ф2���!�K^QB�̉ﰈ��<�7����#��ű�J��C��]�0���:TCTc���
��n]�C,:]ޫe-�!G2z�nS�c�y��1���s�%���ZZ��x[�}v
;X`,n�t�#B.�.�p��3�=D��X\B��5�i �������󬝔�PZ��1��ʊ���"�(�{ŵC�������2j��Bs҈k���'H��9x��R{>z?r ʫ;�Z�F��Y��.}p��%jV��ę �(V��[р.sm���c�ڛ)N,uJ~������0&�o����78Y@^�x^*(�&�?֑��9`E%vUu��ܖ)�m�j��r:���.f���Vh����3z�3��g�<֊�0�{0��u$F{	�D5��DnwM�ȷ� �2�ұ���B2A�<�9���A�?*Tx��7Bf`!	�ӈ�N����M@�I%��	=#�,����̊��\�Y�'��A+�b��U�~NTg���f��-�Q�=W��9�k}���c?����YƎ�+:|�'�mc������s��d6�Fpz|q�2U����u�Ԋ�s�NJ���h##MNh��j�-B��NGC�C.
����j��b�9g�Z�Ć�3��(LB�jzT3��-��F	?�(�3V/S=P?��*Ym�B��e��k�yL�/��c@���g�s���h�!�I��ѮJ��6������