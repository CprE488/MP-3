XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���D�~BDk<����˰�r��.��[�x��J44�i*Z3l�H�7a�ڄ�/��*+�\����RX����c��49�?�k�w
Pf�-�ʰj�)�1-?k��e�
��ho�3a��:�Ì�N�{g@���ɩw��fc���\f�8�h����I��Dw3�QZ!]n�AF�������p��c��ށ;�#Ŷ�mL����l�<�A�^�����ݢMo�)v���@�o);�x�m�E�s	����ӊԅ��J�
��!<Z�
���p�?,2�j�'m,���"�e�mP�Rj�l�ɸ4�o�
�C�Ӭ�(�P������P��iZ�JBh@>�Y�f�����БRK�~���9��P��>�\�-���SbU��no���H��������F���e�\��������"5��~����
%���ʮ�p�_	z7f��Lשa�$er,���N��&�]J4��=�5�	��h���gD�������83K$�7+^G��������ӷ�>\}� {cx��F'�� �w�ʋ&�"��p��;��6�)l��Y�?𭮭o���oJW!cPh��3�4]�����|�����c}�J�#�p= <f�-!��L����+���
�x�hGs�^E���2�S�(.�.,����Y0�fϷ�@�L&��7�$�vN=Cƶ�s��u\�b���&��}Oˎ
ۛ���S�I}��F)R��<'�&
?�RP;���E|0i����	�)��wqT��0|�@D9�ĒC@�H�����O�XlxVHYEB    2b39     b10ͫ��%�T0�R �H2f<�X�!�9i��0��/�D��D��C$6��U�d���9�v��
l6~s�i􋕐0�ʴ�V���W�b�!���~t����G�P��(c
��9rܷ_O��������j�~m5�lf�&1R���e��fm�~mg�
�B�+������F%�lB^$JzLω�� ��v�����?��'�  D�;|4�Ȅ�A]f��Ԡ8��o��V��P*��cPŮmj�8��B�_=sh>>�?�`fC=K�O���ߧ�"����j���$����?�1Z�u�A�^����	��{�M���ǟ�	N�t�qᑿ���!.� ��˼�h��s��Kh�jXU�&��|���>>�ox����'ZpR��~b����q%��P�L�]�y�F���]��7| ���"����7��vV�*�!��<tMC�4�����kWx[`����������n���v���3�Trou�[p���r|�<��>%�{��I����[��X�'Jdg�\��A�E�b���ؙO�zA�II�-daJ����;F�r��.����M]l��Agj� �ݭ�ieز0�<h�VF�8̶�]nm="�cӤ�uX�����LOOZnT�rw{�)�<�۬��5�]��W�Nf���WP�c4�
c.ye�Ӝ#ma��6��]+�.��v'��OPPh��3.3 ���+=n��7Y��]:U�5�>�P����ڨuv�t��Y�'R��^"	��l^N�ŋm��܏1.9��e���2��_d��
W+��
)� ���� �3�k��+��L������f���.������R���
>2)��>f�Blv��_+�|�4�J�|ǭ�N.�F����l��M��	�1�Uf���7:l�N�,��t��ESzP݄�V[n,*��\!��-o#m�|*e�=��A�zq[dv�~M(�3k�ŌPc���-�H
��ԓ|a`xѵ�M�:���*<2kx�<�r '�M?�e��M	�Z&���ų,+�E@�{��l3JaIϨ.�eӟ6��@��R��R���L|Vh�8㓞	����R�2���u$DցyhM{{��	yb �aH��j�H)C"@p_7�
�{+3S�u���'՚�+o�A��$��9z����
����n�.HÌtF��;�U�ޝW���7y�4]�|kH���sXѕD:D�D��Y�6*��aۯ��h:�q�=J �9�p��3���Ai�0T��9ݓ�>�0���m����e�B&�
47f���Sg�q��,XyZ��|w���s�1l�t�`>� �9X�'t(��&!Oa)ȗ1scc����,�~��-���'��j�9�U$�����H��LȠ�bOV�O�a�>'�t��¾��%���~�}���l޳r�V����Zҍli���Ea8s��?��,�,���#�n��.:�*q��b�6�ȟ���n��p@+:BA\�<:���$$�P̭��p�G�h�2�@c�r5��Y��5�O�{���P��dU{G���)��z��K��.�q3G
�`�k��Xk���a���6L	M�@�Z�0��&6��p�N�
�}�k@TN���Ԓ���|K���Ƹj5���&Ľ�E2�EV�E(�e��*���dJ9����1�Y-��o(��_�j�[��T�C�?bB��W�L�BY$�� ��P�A'������	41��?�~����rL�p!��r�����Ewb�ӂ��M��2����MZL=�W>��b�1NCHN�ŝb���dM��)�I�����rHZr���sȦ/Y�� ���h4N������,�)��@��լ>���f�{Żn�g@Qw	�vI3n��7�h�l��G�ޥ�;ni��ﶃ�b�U�@yX��E.x��Y��S-B=�i�l�2 �AOa��h�E0Z��x$�1�j�$�-Q�����@)J0���L�����ת�P+�c~�C/=ܣ�4���^Yj�
÷���$��<�J7K[��
�LM����f���SJ���g��F(5��Np[�CM5�[������H�{��#�����W&��-x�[��W�W���9V �C�]�ڐC�9�f*���}�6n��fE9J(Vɉ��Z��1�U�]�ȵi�6�ر��?=s
���$�U��r1$u�q�8S�lh��~�	���emˡ}��1����֘q��2QGIP�G߆���
h��� �b������pRk�mΒP&�r�-�Q�)iP��B��y�������]�p��v[��y�����2�?��#~�$_T*o�֐�
�ԏ�I�>�[�A9�8i�+U6g�+�8���f���Q��>7�tR	Ƶ{���]��蠟�b,�NbG.����
�z�J츲=�N�fX�ɷ��X��r���X��2<�X�ț�ʋd2�)DYJ���!9��Ō<���O/��@EX`��xM��\�⾶��L��Rp��bˍ��-<�����n|��a�N��\<��$�=��S[LB٦����{�����g�,+�M�1��ǒ�#i\��<�VN��.8�뻔�N�a1���a푣VQ"e��Đ	�
f�v�N���s_.�냢�i/��'>�;N�T�E,H������`yD�rU�]|�J��e#ml����P�5�)�]����.Aˎ�zI��8a��E�06Z�^{���ї8�Dϐ �~���]��O��p��=�^�y�"��>��TwG�L�N�d����2�h�x�bI������7�~1�9?��