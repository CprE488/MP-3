XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$��^��gj�_���[�$>L0.E�c�Sd��q�]�2���#�5�w�v�ϒ�3��e{5��O����A����ў���ߺk@�ӆ��zk��V;A�ДYQ�:�Gi���ՙ���k��$bdv���<�(�h7��q�Iaa�7�\-%�~�ǧ+p�<m�~�r9�(�����'�X���B����n
xYgx�ӯ��8�B�\�Ϩ��"��_��"wϰ���)8N�ZX��4�dC%�~4�G@+�+ln~8P�K��"�AMAHB��8}+� 	���-e��O2�����hK�N�:�i�����MB	��)��2�ISc\�����,u�Tj좘�\��#t2Hs���7���@�aMpB��6w�ӯp
��)�œ{�q��x�C_�:��}/�2�M�O2�����-1��� ����ԅ�B"B����}�~Q�k,�����<�
?�''9�*�	]�S�Wg�~�AӸ�� �Bqj<\6{z�Z<�v�S;��Q\-DR}����/$�	b�"�*�_�29=�,���aT��:e�bY^��n,xI�D�t�P��Aw����fk�'��Yh�a�i���xoB�a�0�Iʽ�lӧ��t"����v!�4�i1��Ľ��,j%�"T���ƋA~�Js�"�<"�3��0�$�iɀGoMUGES�Q#�Z1�E^á�U����T���]S/�^���y�bW�[ �R�(����e=\�����~������PO�ٛx�������Q���XlxVHYEB    5d54    14e0���GZ�X.w�a���[s�r��B�w�OQ��h��FL�7v������:F0ӡ%s��c�B��=�@^0�f�9��&1'A�k4l4���&[5��4�ޥ!��%t3MY֎� ^lh+#�<�`y���ٞb�lp�1.���Ǎ[�]��<���cZ疝9�By�ͽ����IN��zV�ZUiA2í�����ʝ���J7���v�����w57�Y��E:��������a j��@Y�poi��R��Utנ��Z�s����Y����ZMBx�*#�	-�!P-����S����G����>��g9v�dR��u�s��ΟQ ����AD^���_�f@ܪB�0�Bxr��d`Ʃt��Rb��W2s���
9���V,��x�,U%�O��?�����;o���<Fc��k�ۦ�%�[��b����WsM�K?�7���I����6��I�Rߋ�^7�����?8I
�ۂ�q P%쪘���,����	�u_��;6e7�Dz�M�4?��R�	{/�F���<��>q*�Ӧ���
 ��# �9��P��!f��,���W�� Tb2�g���1���#�X��W��X
B1Œ�Ź�.1�����c�{��Q���>t�L���B����L�tS%�dP"lu��V�P��K��E_��c�cEY:~�GN�f����l@��-��@CЅ{��,���~�x QO���<H�ZT��l��D���3���+X>(A�]��xρ�Hh���gq��ᐅ�Ń@�/�9p�X8I�|�ߦ�f�#�ͮ0��@-u��N���TB��Pf��`Vsz�d8/���w���PK_�lVCUR;�qW�G�͓[�b�ck��m-�����_�����I`�^eTPi?��rcH^��;x-��@_4毈<�����I�VF)\F�r���4=�J��v�i�=�M頱���V
lD`����􈈚F[�}�������GC�v���o(�}P��+v2p�+��c�#-e�;�eis�w��:�UYa��P��F����V�P,���V��z��E,:T�^$Nd��I�2�؈P��� +G�*
%�ã1y���?��0^��pl���P1�Vl$p���Vz��mD&�����{��m��ߣ��w}G�9|όb�|���5FG+_f_#��`�K¼:�x*�6*���o���孋�y_r]�N,��j�aY��v�6�ZCs.�!�d�p�د��N���'!��CАl���l�� s�Y�1���W�>}��֖B�$nwt7��,��ln�ll�_Օ��$�����iW%y���]C��{~ik 
]B�o�������^Z�R�����lzF
���'���K&�w��|�ݘ�?V���*R?!�Ave��Z(3�BE�l8�&S7K��+��&�c+><'`�A�	����;
>���&��4a�ӿ����3�ta�w-J����^dt4W�w�C����6�hX}��d�{�s���FEj�i�����f�XVJ�g��O�^�AxM
�K-'�9���%�,��
�F���Xg}י9~O$��V��4b����xhf!�Ta�*��:/T��;�1�G,�p��$"�TλC�ZJ��zK��O����
�"���(�^��5Sw�/u�I'C����Z���Y�t%-��T����� ��֚5�}�2'����y<��_6��Kc�7��z~;��G��_.���� i��s�Go��OJk:�$ŀ�E����d7�J>�˩���2Q�}���&N�l����X���AX���Lp�!��춣3ױ;6��j>b\i�Y�_�ux�ۚ�(���̶q�*�\�2,E�����)2�XbP�8<�Z��h%R�Y(KТ���!{��䓭���1��vt�(/�¿�^O��TF�]eZl�IM̼u��Y��0A
:��=�(�X����B�<~;6�k�!g]�vi��V`]�P�r���l���,r�h�|a��Y�#�=�9(-���{/ఎg[�x^��0r�+�����|һ~����*�6�.�7���V"�������TR��.�l���d��f�F{.qpd!J�j
�n�	��J7Bq�#�Z!͛}M��-�;�-��j��	���2�X^w���$��q~HY��T0���`�
��� �"����Z;E� /@`Ӽ݈�J@gK=�bcj�/�)7\��g����gv����LN���6����:� ��o㢔��h����nF���YB�^��Q����K�����P�!;C�}v���M8舢wݽ�ݸ�8�B.�<ܹ��P��m샂��*�96釋rǉ5�7~�m�گ�q��o�Bix��2�i�lfdj24� ��/��	�y�E�Ъ�h] ]�r�6:�&��Md"�c�Tl��9����h�\��
�$����xxK�>�j�xڪy�
�.v�7Al.l��yqRͱX������_��}xp8ec�
�<՝ﵸ!_�X��k���@���c��X�B)2�*���8w�O3x����ф(��~�A���E7�!�E��6;[�HY?惣���u@0��5��齷�ޅy�Ǽ��&�ƣ'4n��)��hf�	�o,���ֹ9<E�θ��%kQ�ȩ�mS�ڲ-�?�j:C��݌��F$�/�r�s����e��=��b��vU�u����:(�?23��WS1�8�
����&��Q2ˆLÕV���3�Z�E�	�@�)D�HT-��7:�\E��Or�����S��Ӑ��k���#�Te=<��Zo�?�5ї�"6$]����-8l����QF�]�v��cs����结;���9%�G_�4͎���$�ɲ�U58I��h&)q��m�p~�a���kx�:3B[�T��4��DC����_��M�y�Hs�F��.�fݪَ���.���Q�Q�yfͷ���#�d �5�Os��M+����)�n|�y�Iwʼ��e����3���\D��-���;�y�X���I�cȘv|E�f��2�|�Ȁ�vK��'5�PX��3�/��F��O��yOy�Đ�z�S0G����Bl)O�a���BH�1����P ��$����i��L��a�Y*��U-�Y��VrM�d��l��}S�>�����ؗ�+����?V4�D0�O�a+>f���E:�V#��T^Dsa>�n3�ߴL Wv�^��5e)K^�y����U��g��,�xGZ���S*��ٍFZ	b�ZM<��*r��ނ�__h��9��{| MR�\F��[�tk����<�%C�U)��[�U7�9�][`�H��UK�i
��h��@�ߏ�����1��Ç&���9cz- ku��#k�r����:b&I^��Y���{��8ޕ�9�y�}��_�I�BP��i1�Qe����3c��Y��n�X<]��pP�x����ߜ2����1�6���j~��-�^8�nN��l�0� �	�@r�r�:�d�W9���]���_��Ή]oJ{�?�}�`�یѶw�;Q�1F[p�^�!�p�䥓(_"ո�HI��P�r�i�d	)۪H�Kk/F� ?�cya�]�lz��[- ؁O{�7p`����=���l۾�k��fB3��sݨ
��Eϫ?�3���Jn��"��H�����(Z�,�-+'H=Ϫ�a�﯈�ǖ,a�g��|��)�xJG�#:�"�Ys:�wyR��eQ8i\y^�������yX������u�I����$LV?��2&������t�In�t]��E�|i�/�<�������R�e�-sARy��"֎A��Ш4�s�=�� b�_��^$q,�z���J����>�kD�%��A�N6V����*��@|j�h\���?�4Vv*#f�^� 'D��xTñV�d��C@$NG:{֨�Zƌ6�i+�D�m_����F\n�����:����j�Ű��� �\U ��Aމ�Iy�жZX@��Uj�|�#ʒ.�Gi��f���s�^���i[!����-L�*,0�;-�}��?�O�`ts�'��r��"��d�y,S�%�%V�Yt�P���6t)�&N��"*M�knLq�9!m���@�+̅1"�v������}�%Y��0�6L�J#s`���&5��BYg
�����\l�Y=������:MGe��(��de�
���8+*Mb
	�#��5M�~�����wm�5�����pid��
��a�N��0:�G�yL�]�*�I�w������Vs��#�(9n�+ }fE�v�d���'��h�a(Q�y`�-:�������n?��L%C�D�sE`*�<ΰo�.�i��
~6ڽ�\/�K粗v�~��2�a]Dc+PV��(*��6ޕ����	�~|��m,�����СH[޸��ցO�U���$�v��:$�z�����}U�������(q��C��-��X�9&[(��CW�����Cq /Q�a� �,y�;>U9V�D��k�܋v��<��Ŋ��uQ����*W�σ'O5>�ŀ�q v�%�9s�x8��g�	����-1˯�}U�420�nXX0H�T�VR���X�2Td ?�*���O|���e�ݭ�ͫ'���SE�N�d� �Y��%���B� ���IX���?E��w�=��X��CJ���g蔟�뭿M5C�Y��r0~�i���� �'c����-�I<��KPi������q�<Sc��u�)�]I�V��m��:����.Ї R1����o���<��:�ގA�k�����|�N���>�
o佼�-$�ux&��n�j@����W�r��MjwG^l7p��/�kh���JlաY/0��D�a����_�I ��Q2�ׇ����1�(Ia�C*���t�h,fz�xc�l*7�$ZN�^>�8��c�-	�1[�T������H e��(���R{�k���Vmmv�d�N����:O��ȑ�Q֜���TAh�L�>rdO�e���<�]��x�87�����G��`�����dcG�[�z�/�m�W�K���!�D�$����|��D����͊����>5�e�@B0EU�N��2��(�x�DU�ź�>��g��S�9'�f��h�N����@/w?�0£J��
U�i%�IqA��#	�t��ps���Q����4�Gn�kƻ3��X��bV�f��ǨTT�FaNݨ�Z/�)�..���/҇�W�e�B�̈́��}�äx��7��
p�%�m