XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������|hz��7DOE}_���Z�k�h���~ݿ��������([���:?3�2d����i�jY��4�wl�l�*��v[�O�7B��Ji�FEi�":��p)u���NZ�\��LW��l��\4�/���>k�T���ª���Q�{l⼯6�{?�-�ߨ�uCJ'���ԗ� ����m���������25�IDݗ�<����5�%���)�b2�	�N��{Wf6@�ߠ�1y]����z�39�<�0ʬ?��N�L�����1T�w�׼+S�sD+��E=..彩��(�^!;�"zGf��I���20��mP�W�I����:6���8�T��v�@��>T��u��kU5��ob���Q n
�@�:L�|�$�5.w_�*���m���:��O8�P5�ɚV_��N�����_�7i6^7_T��dѡ�̕�,���j��	��D~���agv��se�5�X=e|q\0�$���n/�FJ�
���v`26�6g����"���p|$��C{hy2\��Z�*]��#u��C[h�tw5S��lЌs�~e(�R=�*�7���ל2���t��,_dmxhT�V������U�����he��_ٺQН���z���L����W#6��뾄�ꎵ�_����&���p�%��?s�����ə���OӤ9�����^o5ا���1�Q)����J]�D��q>�1���O�{3}�QrX� �-q6h^E�E{��8|vW"�d��*`6`{��+�)XlxVHYEB    4b7d    1310�Q�z)��N��p��#;e�N����ӅӺB^/6��@#�4��C��7,���6�}GC�R�L���Κ離P|�^�t�9'�p��_�J�W!��J���9X� ���#�Bӎl����Q1='�"O�K����a�9S$.�Ď��n��ڟ�zjh|�&�:Y*ͻ�ש�Nr��j��Y��z��;z�<��̈��9��Y�����z�	���5ȼ򢛡8 T�Y%����":\5���Ű������XK�Ѫ���L��C��+\l��=Nt�K�/��au'�;���a�s��E�bl��Z�';��i���8�&:�4�e��'1�� ��8gS�Ɵ�Ɣ��ݺ��o]s%w��1Ÿ�5��t�`a��,��Qr
 ��W����F�S����X� \$B���D�S���0؞�����PIp��87WR����/�X��("E	��a���"[�u $��oV'�Z��A�+�՟�ǀ�#�!d/�1�f�%t�[��* U�B�l�A���$��+�8��Z���\4M�$�Ngҭ�//,h�	��硕��5��(��p���>����5Z�ɿ�����J^h�����gϾ����C�b4���m�T�~�G�2PY'{��]M�fr�MO �k���}z_��d���������K���h�ց�&x?��G�rL�$�pvg��*zO�6y��oe�?�����F� ����R�)!
�-�ϲ5g?BӴf�]��sg���9����<{@c����(I�4�.�=�Q��K�G�WDD�H��X)�ߓca*�w9F��6��{Q9�L�zG�b��U�c���"�s��GF�o������������e�L�]Z��u'�I���rC+}����B�w�^��͍�1b ���n��<C۠=6h��wK�υC��%F����BG�J�I�2A[ن=�8����9���7I�kE�y��n��3�Q�<��>�u5az��%#�G�W
q.�`�>�r@�g7�p�
���E?H�YUq�q.�����uĺ4��)\��N��'I�e� m,Q
��yn�@�Y�5D��<�T��gq+;��@nO�^eL)hm7��C�c��X�f˾�����3��tKqX���_B9P�3�"���C�A�c�	��fj2F�G�)"r]�I�����2��uf�AC��!����T�3����oƐ�;�*s�[�J��R�	M����k#�>g�9�q�Y{-�E���q�����x�9���[.��2��OI�	`xM	D�ǉ�I��l	�$�^����o&:����G�����l���)��Kz���������Ҫ0����" �$8�z%A�[�v�i��o�����~dY���NN�X)ٟZ�C�|Z��|= D_{c;�-�{��$��+�'�S���9\/;��5��ԓr8�I��׼rc�}T|f#]]zNCF�k�DO�VzY��k�������uՒ�9�DiN���/7�x��
�O��~�������v���@Qt{�x:�����p�L��l�U"�ކO��ߨ�e��d"9Ψ�Q)�i�m��ǲ2QD`\��Os^���f��^�����iB�o�F�_��keu&�T�Z�Pz���z�^͢���qf����b��][��![zI���I��s �D�|8�,!T�Y��k���Jr;�c�( ���0��F,�����֋��b��E�9R�"�<Էz/Xf����r���L�V����9,�Sb�jFol��r�^�y�Ј�f<'N;�Z͝�6�t������~uUTtx��US���CӞX�>о��퀤��-��NO n'ړmC/4 @L��s�yL��9��5�#�鋮��C��	� mH̉G,�o��2p�h)�?��%���S�*y��kO��lDf����L4�9��`(RuMH-X[�CGP/p��\~��}$���t!�����C���F��Ì���^��#3�cP˞$m ���\��JI��i�g�[2e����a� w��h������
h���$S��r�/E�#&�Q� �A��o�Q=�Q�$�Q���1(Y����1)|U�T�LH���v&��a��a�)[�cکVI�ŵ�t�^]��QJ����H���]w��,����iŉ�=�He�k��n��PHj�<�6�:��y�a������\Pq�	9�tǘ�|#�TQ_��p���ܖ����XqV#��v��)��w�h*�3Jib��|�<u�L1L���3rc´9�|TX�����q��]	��`��*�d�R�'r4�ņ�G �������F΃��h���Z�04��	�C8��^�h��U��oh�Op�
���z�^��A�ޟ�=��;�Z�����'G=Y�]�5$�!�=c�j�z_OE7@���Y5u�&HN0�����e�(�Ąȁ�j��`���`�Y��"����g�����/l��3ڀ������
�2~�v/��g^[�o~`�~}>�ѻ�m��8,�R���g+��V���۸��a<��)��8�LO��`,�QkK>��G�^�Z��y�i�	qM��0ǸϠ�����F���B��ó~34�� �f�T�T,��1;N���(�W��gl�X��+�m�ؘ3�`э:�d��o����Gp{�5lR��3�(51���z켗�q(?4���z:�`z�w~�������M��p�_q�@� �������h[�Ͻ�]$5���s_��`LH��w�ѽυ=J�Ynؕ� ;+x�H9z߃�%I�t̓C���}��q��4,��}�;1�S7�"��l�w ��b�� ] ���>1�!��XܽLH�M�qS�.(�N��^x��dɼE��AW�Iz�!�q��*��*�U86:��9�9�٧�,]o;Cjmm��k���U��>��m���|���`G@9��q��ۭ��4�����Q���y��� �M2ғ�� �y�XZ�*�F��a�݇P-�a���:�̈�18�1V��/抓o`�Fj�Z@&+�Q-*�݁
3ݙ"?b�
M���˶�T�'^��U�hg+�4ǀ��ݽ�*��y�B�"u\iT]Y'��JލW(?yID3^��3W�;W?T�%t�s���ťׅQ~t[���`"%ղDӓNl#�y�z�͘-A�����R��y߉���Z2*�TZ��L�w��o׏12��&�x�{�� !z'�٭��@�Rl����I�P�Y�~`��05k���x�=IR7�C��,�J��^�^��Sb�ma�Hm6�p�lg�!o�:�z�9����� T���~_�����Ify�g`�i�@8뾓c��� &���Yz�\X��&F��"�� �T���J] ��p�Z�ciF�G������}w��ZS���XT�6m�<4�mX^𖐡���@��tО*�T�}��&��QX�Aa�ǯ�3�_�hUF��r���>-Gf̏��Z�]�|���zL��N�lF����w7:~UB��>���kb��f������A�YL�T��w~�"�g���TP2Z�̴)��b2�]����^ֆ|��V�C.M�IV�J|yC�VM��<�#q���X1S�aP|� �h���%�����+��3��3��4멑���l�߯����l������4�JK�߸Fr)z�1�����G��>������?�Fe$'���M<4�.ǭFG�*d�Co��u5�
5	s>�Ԩ"���޺:>��у�K4�hx��l��W���g���;��*dV]#�p#�Q��A��!��C�Z�����@z�h,�L7R (gX�J�������\0����Ӗ���-��^N�3�6BĬj�!�����K1�eT�~�A
� 1�V/�B's��tH�e�1��&_�H���=�q/��ޱ�ĳ�t	�QP����B�}G�%�&
F���~�Hf��>}2��!�����%X�9����4ba�g�Q�/�q��� �(�
�0�Z�P��ҿ��W�j>���;qI��a�=�_�)L���3��ɏ���z��>6�ΆeJ���������XF�ng��#�{�>�
�e~P5��3C�݊m��M9bTVuh�Ɂ;���i�h^�#���{)�>��qnxcO-����&N��I��c?Lٟf��Ū��0������iJ9����u�3��\??P���y�������E���"M�WT��t���H�Tr��fK�D���C�,�O(P��QQ�5�T}�VyД��W>n	E\VQ���,��n�O��Q]*��U�ݯ�o�G%��Aէ-��6��\��E
]�KD;ꃌ�s�v���&g{�y�n]�1-��O����q��� �d׈�8��L
�#Ց`��!SۯX�{�:O�t��"�q_��o߯�`^�b��-�Q��7f�ճQ9���K��~7�s5T���>�1L���~��% ���L�&��
%���} ��w%�\ǖ��8�$�'$�/!�r�
c�&THl
G�!Ȝ����"}���\�^rTKn;���}�z��%Q}*�l���ڵk�� TE��y���᠋c7?��	<uB�~�i��r,0����R�+8���a�Ԋ�9��3;;\ۡk�J�&���^?�³]��2@�{n�ޑx����!�)�6Y��'P�m�ʉj�3���'��&*���
Ʊ���p���z�����;��ن�D�U��"8���TW����V��\f�i�[��ب��]���1�&s��o�f E驯�&*7�&"y�ߠRo�&Ȼk_	�z��G��l��O8c/�	s��N�Ե�8�M����5�