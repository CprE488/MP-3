XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i��./���>�m�������P���o�!��� F�);E�
��-|�v4��iyN�}
�0	��4���\�`���If���q�eyi:�hwh�Õo���>��69'h���> 8����n�uB�ֻ���c���ןm��}����{���HU�y��(.�: �գ�F��:�BZ���qd|�Ď�IZzW�D*)e��nčN������Os�B:�
Cu�-��v _`i���_�wD�t��h2��b���|��:I��988~��-5���fl#%��# ��,yꢝ!-���Q~�Eh��w�����s��N	&�bfF� ֩�U�5d8�Z��g9��P��Jv������, <P�oK��L�#B�+"�;� �H8�Հs�ZC�E�a�Qf�Yd�+�.7�m�·�[��2���2g�2͜��(��f;'.�Pjw��B�j�ḅ��W4(�e<�~��>�#�w滻�/����ރd�m��T�%��D��Ν��L�Jj�V���)q�Ȉ:�����]W���p�b��r9��#���Y��Ew���Z��]k�ŧ8�6P�(�;��T�qM�j�9�t>��.���VW�� �T�lH	�xz�}��"�>�-޲D�@M{w<���;�!�e�H9g&߂v?���B�g*
6��ϭ~�u��gm+5EJC,񨡮ߋO�?/r��)ZP��(����u)�1̔t=�wR��ϑ���1c�JBZcwJL˔�Tx�X(���MM̟7O����{��S��4�V;,e�ԎXlxVHYEB    48e3     e00��*�z�|-��Be��7�#���R3E� ~���0;��H�dNT���\� �l\����a��[G�v�Zݼ\��ȅ�ګ\��y hkE��:�&<n'z�4�N)3�ütRo��Zf��LwtѴ�"�#�XU'^&]�f�4x����gg�*�cx3�ul�H,�6i�@�R�1Cτd��}K7�'������m��U4��_��F�������mCf��XŦ���8�ٛF�[�A8���]k�j�,�}��f��iy�3�d��ePc����z���ւ�mK�7��0 ���)T��{+��e��[�J/�����b�^Muj(���2���_)9�M9��Ewڮ���M��{�V�׮���#K�ÄV;P�0�������mw~q>�ǮM_St'�Y��V�a���ϥ\���ɦ��ѿ���?��9�f��'H�[�z�����w�,t��m�����ӫ]ث�T���0�u_� Y��[̦z�<�N���V�/�c�C=�9#���d�䬞Ϫf�__Q�,����Yi���'6z6]b�D����4]�9J>��6A�8����I2��1��4X��q�I❯OG��G��/����EGL�y���kQ��AB��ma]Z�5�c��m��)e��!d�����G�����'BmlC�'Q�_*� ���U�osX�=��78�*�Un ��d��M���3}��F�<X(Mϙ�?&ai!��!��jQ�|B���Gc�1U�d�eXsJ{��:�m�!�f���MV(�b8�l���Y�c�����Zyz� �F����p�xeVv:���O¡��&�W����ڢM0&���U���������>����f$CP5�}��o�},bi�ݠ��:�hDU카�5��s&H=o��gT�_$���f����x��:k�'�=(�L"�2��Y��\�Y�iP��C���ɜb[9��V��;���Q]���/����~V�۪fG�r@m``���U7|[B0~�_��M&3�\�����`�c̟M��E��'��s��L���� k(Tk*��������q1�н~ԟ��F׏7��]r��Bsw�T&���y��%I]_C����2a��X�KΚ�0�d �3G	LN�_�D�ƿ? Kq�됽�-������5AY4��\�ʽ,[�<�gA~���]�uk4�!1i������=��ҏ�伌����y	�x�|���Mb50�^J/b70�:��QC��b�����S���gn�EN5 pf�"�{^q��ڽ��|is
[�d���8%���]���m��wRv���`yik���p��i�h�3��"_'�V���+d��zЉHﾧ�`;�]��F�����z����>wkC��2/9)��'E�����j�@D�t�y��*�K�Z����}��$��LNxԋ�K�d�g�.��d�8�uz���n�����tJ��Y�u�Ϻv�_�%�D;�����m%7�<ă��M�68#ީ��홟�,ᡟ� ��Ï/iDO|��7��j c���%��3�d&P�BY��r�e�j)*^~�F�s��+��A321ZIJ��_�?������{/�ʌ��x,r�4��@�b�3��WDͮ��D�(T�僛G'���[�6�����H4�s��r�.���u��z�H
[
��m�8����K��7��4�����N�Y�^YH���X�G�_TN�CQ����T�T}nx�(�b�kɋnԜ�N�2,8�>L�/x�2���H���� �Zy�Ո���O(��`���H���[{�*2㴄#D.�y�V����
ב���bK�6���
_�Ѿ ��R��2�]?i���[s��8�:���/�����PO�������F�'3V�i��	��2=~I�ya�J��z�����f�1���e�|ԡ�<$�I�E�.���V�%0_@�:%9���h�����9k�|Y ��Ȕ=g_��)~�P���Y����S�I���jW�Z?0h�z���.��O��{���N.F��Yw�#������.�.34��a��_?�ډ��t�z)�!r�O����д��W���9��i��5q݌�s~��?XS-S��*UY��_8jo�yiAa�c��p�*��P��'�n�gy�Y�rR�C~<8�Oo+?�a c�+
Əj,��TF��T\Յ@g�n�Fؽzu
���+h�.y?��	�A@�ۣ��G%1���� �u�70��)���G�*cP�lҠM��#����aI@��������1���I���F��g�Ҽ�dp����j�����U�q�WfpG�o3Ř8x�\�OV�����SF��c��5����o�����c�g�,w����|(NCQ�*Л{)~s�M@���fh���򀐑��f�r-_2��7���oOeud�jgˏ�ZX�1bDD��(4.x
f����|�~��Bam_�.�2q�u�d��KeD��V+BVKv?\�,��BC�6�pC���0Y�C�Q��z:Q�iuܓڮ����#�]:�����=ΛA� �O?��i|W?$U%����D�i����x�t��V�o.����߭o�	����$��t�6r�5����̙0���y�N�Q�aQtH��o�V�E�'�P�V:D�*��\�=�;D|�!HcFu
`��A§��|w�T�`���f��~�J#n���4�]�荇��(�b�B�{�BAѯ4���fw::
��eI�}�e�=��9��!������f&�/iMD���~v�QUA_�ç�v.���N�f��2y%!�&�!m�����v�o%E�����q�����m���`ϥ�����������A~vh���}�����Ghf8y��WZ[x��ԭ�^aٿ3��u�����ߩ�Vhz���Ij�SnB����|��!ɧqЭt9���k;��f��U�Bm3a�.~g�(�<����$,ר Oo�DtӍ2kz�2y!�{�, 萁F�Z[{=xA��$���C���O�iI���B���ἢ$$X�����|���8*9�M�����n�Ҿ�=xX�p�0�~?�Y%T7�=K��$+��X�Q}o3���6tU�zw�Ǭ-�R��� ���́��#�E��0a�KGF�~J��T	��D���y������ȅ�EE�/��X{Gn	9w(�S�TSH�:V�9��^ r�Ep�
���ܡu�W�����������<���gе4N��7��_m���+�[l�zku�����m�6��m�}O���+���4�da��e�}�]��z����ie���1� ������.��{(�O<�x6
��d�O=�B��<�`�.UBnv�:��� ɲJ;�eC^m���Y���{".~OD��ء�F��1Xp���MLy����K\RҤj�^�(`퍮"9<;�xʂ�΀wY��'�i�����:���n���K2͌�`�Od�f�Pp�G �	���Ns�#|�3?�{l�zs�A)���RKKk��P�x�