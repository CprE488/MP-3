XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��x¶��~_�v��t`��Ѝx�QW9�ΏX��:�.1ge��D���t�0����#�(�{C��|Y����T�I����o�{k��Bq1��e���q�ˑP:���G��w���M,
��u�o�)lO��(?3�� \{6�M�/6�,�X(Z��f_���d�M�\�{����nİ���R��u- �R�����'o$eN��K
*[��&"�3����"$�ΰ�a�:��c�����n�[��>RPЅ]t�J�p׺�Kק�,��7�Z�&-cf�ۥ4I<d�B!K��6[��d]�_�i\)�Fo�Ւ��NC0wW�����E�A��Qm�ET9�����x��s~ؚ�o쉎��33���Ȟ���e�e��Dob��$��R�t�D��d�[��F<�|����l����(E:q�mLh��/M�px��@ޱG�p���fd56Z�"v3*#VG��WhƩ�Wκ�dKML���}j�_PWR����&BJ:?1��������uB#cU13c���k�����DO �uWb�>�П�%TFL�-wV��f��~�f�3�V��A�PA��ҿ��x��`�Z�"�V�x��F?г�Kɬ�~|�<5�t����������'��"��I�?�;ó'�����d^��Cak��]��&��)ո�u���ں�S-աۺ�%$���L���<����;�Q5�e���L�l$��N���io��� @�<�3갛z�Z~�Q����/���.]XlxVHYEB    5d54    14e0�ꌌ)�<���&��6^���A]83.d\��XGؙU�Y�N��&�_�B��ܝZ���t[���9_��`�zGG���(6u\i��r;��?^na��s������~���q3Ŷ��h�z��B�~�T/H�A&\A�53�I�1�+����=���]�3Q֡A"�@�ȫ��r��Bв6�#LUB��U�\�
u9�����7L��U�/���\��v!�A����׍ּ` �)�^�����ƈ�!{�U���Ϩw��;�*�Ԅ�hD�I�PAaF��b�?_���ܗ&$5� .e�x�>�&����>��	.�5 d�|˴Q���ν�M��/J���t0�M�Z�ȋ��d�ޚ�����|���p�
_�!��B"M&g՝���֧�H�ɐ�ڬ¬�ƈ�r��W���hf��}O�HU�^;/�7���:�M��m�D"6�1X�Ͷ�s���OE�<����[{ǜ�����̿%X4���%4��_ 44����<T�^�Bd�����D4�j����0:i�z�=J�Y���D*aj�~���=�����&i;ۄ���J\*�	|��ؿ�nu�Xj�s���2�����ݺ���3�nlO�m}$�ת*.�`������w��z�� �����|���_�~>Re"���v3�/~
c�Om�MN���y�K�gH�u����2&�%M�]&[���#g���)3iv��O��Ka�="���%'�,�?�u���զ��}��4�,�̯�<D�x�G?�y]���B�]�%�0Hp���_���+h7O��1�I���LbD$�B6�L��q�.�n@R���ڔ ��e6�E:"��q�{�B�E[$:��!��|<ѵxvbYb3�^�7���� K���:Yn��i�G,{N7� ]6�c7V�r���bOH��Y1{Jcf���%L�Ф#=��p�� =a�������N_"��L0�4V�Et���6�`���C�ׇ�pTuy��Y��A��[��j�%�q݁I1���[r޳��)�
D���O�:<~�4r�`J-�
5��xaq�ĥ{��:O}�>L�i%�&������P��GqP���r��ޖ2hwP4jC���F�.�$E��8���y����hP5��y��0�Uw`��P\7���c�}MK��>��k��䃻�ѣ썗� �fs�5#!+�YP���S[`I@L�0���m����ΐ�&����q��KA��)٥��=�zr.�Pm�&����%"s��͞�:��b�n��Ě���(^�Z���9�H^�?�K?ϸ���P�
��$ۆ���t����;�����w��;���V�@�u�4XyrW�ҏ��r��ȯ�\����j�
�k>6�k%��&
C`lL���6e��{��v_��i��0�$�eH�af!D��R��9�ZJ� .����Z���;�3�'�OA;s��q>c�-"��E`�x����`F-���.����H�_���m��*�aeW?*Eƙ̯5������,��2��)�(D�L�|Nv��x�$�못:��V��e��j�~�T#�+�����H:��<��ϲ�Fy�ȳߒoo&w�Jv��a��U����`{���o!�[K�\5����Hi�z@՘�Ė?����U9y�hܦ�	���Z�t��&���_�Vq-I���9��ǃ�;�loٸ&ȤkQ�͢�g�|���l���`@�y�ذ&k2�#R��t@mk8O����ŉ�z�*RbL���3nq2f�S&v�m������:�,�ux�;b�uVE�����G�φ��Y���ҷ�\<6e�CȀ���::��In��q���#��i�
;�E��p����������ޛ&t��KH���Ó��+QX�a�WFF�9���@(���g��?������:_j��I"��v��������(&���sIPM�wS}+�хI�n?���M�J	��gely����� X�v�^��/����Z���݅���+^_�`��WqG2�������s��s�-�E[�1s��o�\YP�:������G�%� V@�Q=޳,el�x}�a�C}�����WX�X�@.�7;E�`�fެ����C#��mz�z1mR����t�g�ޢ�א3�x�2s(�ڞ1��3j?=D��A��s�m���@6�������E��\ׇrYf$gzt�Қس�dj6��|��6P[^>�pZppb��=��b
��N�_=Q��GT����D:H�jUਭ�l@�δF?�'@e�)��&tm�:7N�g�#��R�y�&R
>�Q����*�Z:���#b�6�#$�$���U�Ց��N���̳륚�=�(qH�%�͗H�h�d�˩u~��?H�V��TX�R�:<���?�+i�jY��@�XNΣ+��_�b@g=�01�A��J�����O��eW�e��-��8��R1��M`����N��)�ff=�m�ph֬t���5�_�������_���g:I������S��/;ϟD�8t�2���*��M+�<�������[��lR)������	����$C���a�K\��|e�w^����^�_e�u�q{�/��vyh.@��'#���⹾���i�+�e���v9�֥n�ҷ-�Gn�߃�����<W��"Y�ˀ�X��br�e�}�3�	�-`Iq����3x�'�m4"�cB	�ڔ35�;���6���.��G��}6��!b�(D����,A�ك�DTՈ��xq�Վ�C�pߦ!�04e	�;ݩ�ȯ�E�U���`jچ�A��N֌@�aɽcJ#�K�������{c�4��+�nV�(��H��̣�����l�_嬢ʯh�Z�'��q.z��>	:F����c���R�Z��8��:�4%���ӽ��BiI��M���4�pӆ���.9���ԩp_�����Bz�@�����|f��[��o����] 6�wW��ݒU6��WX�T���c�Ұ��z3W��`���5�:�d
R\߭#�&R���|�#���a�C���W�f�U߯G��C�e'����c^����2e(�8W��z���� =º';!i$�$�[k�j>%P�5����҄���h�����h(ct��� nk[C��:2X��q@x5���	�R0�<�d��m�?u�{��Ȼ�u_ΥB��e��;r?���ʰ�f�$b��vm�L�y3%��c�$7�.teW짓���s�	2edJ�nQ1�h��>W��r<�!j���<���/=A�}���qN�U�O	ç��~wz�ms�8W��7���b������=���}��vC�M��"��
�i�c�ջ����ũ]ŀ~�H��`3���cc��M�d��?&*,�����1Ƿl	p)��ń[t۴���a��A�H��(���$�Q�7��f�Z��Q\#KMy��5��l.�$%�ֻ�)ZQ�P΄5�,���M֊db�Mn\mqLmAl�3Y��̟��kN�ռ�t�������00�LZ�j�L�w���E�vvY-�{�볚�(1tE�����U'����H�T������-ߴ�iaJ��C��m�1�i�=}¿���]�����8��F�Z������[���n�N�p����Ax|o�݄��J�$X�_�|a����ힺjd6'�>FՓ&!&|O��l��Z�~���3k��Z���D� ��0��bՂ�{+O�O�����M�K�~��m��� �:v<�Ks�`�nV�f��K�q1eRA�Gx�	����L�Z0���0p��Oww�����K,�����O}�RG��j�np]�l�!V�!��|C��I?կK^9	�1͌[o��8�M@��W�䞫A<�Ȉ���6����e�-Gv�|)�YK�C;�S�հ�4�IH�xдv���[�^#4r�8M�Zx_[�!���F�+�L���c��He�&���<����	��8C*���+qY��~J���._�]�(Q9#�4⤒�]��近p1���9������9�T��f�F!2{�Unb�L�.�����	���o��ᰔu4�ݱ}��g�~� A;���P8p�{��C�|�K�)���ݙb7�$x�����Zso_�fǦ�Av՞J]�˸��1��ܲ���%�����F�J�pk�D��a�o	���_�)��cӠ�����&�E1}�`:�%B��e �i�[y��(;�>;��(�L%���9����]�?���e��#5C�N��� gթ�\Ȏ%Ө�p�߇�8[AaC�m����4F�|�g�fdg���wKG ���V��4N|���`(b��2졳l5�R8p��纜�tJ��6dT5�
����2
�m����!�~[{���y�i�yD��3t
��76k3x� �����,��ٲ�]��Am���U�
)�{�c�\6�����kލg܍�1g��6��㑙{|W�G�Rך{l��#ez1SY�:}8�����\,��q�e��~����n������I�|C?��l�L@���������*H���᠁�B�f "��j���*Q�%˚Ws�)�vޒ������G��W ��Z���<��ҡ�ej�[��u�J[���F/+�M�]��-,�+d�t��\�0��M�����Q���[�"�߀܄��VLtHQ!�#�o��?��tҶpɭ3G2)4�S�6Y^�uD3e�;\-��I�|�R�D~�����i6�:��g~�(^��K�������t�saa����c.#'@�ޔ\�Jg���LLwxg,I,a�@RY�,?Î6��`w�v6a�3Ջ�h��y�P���n�{��WόIQ�xSF�9���~"�V0Tnqç��|c=�#q$sGZ�2�L����ɍz��S���֑p���[ՀzYq<F��ݤ�?�$�"+CϾ[Xp~�l��ó��:'o����bi�����܈�Ų��z]E��"�',��|鎙�㸁w*E�Q�5{��BۣL³Ob<o�)岕�;W!VM9�2�����h�5O��ɡ�b�"�ג���XX#!c�F(��aw��egI�ϣ�z�׷�>��=��k�W�>�\�@2:�KI����	d���D:g(ǿ0>����T;�
�<v�x���p.�t6�?q��x�."�E(����n�!b���{7H�f!Ԥ������J�z���/�R�/�7�ѣ�w����[K��&�Vnŀ