XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A���#�,(�`A�~��`T(�j�z-�L�L ������Jt#�r�L�0a��!�m+��0�E(ru�*E+";I�h�)��ʙ�O����2GG����-�	�k��-�7���+N��Ne����L���n�OP�7x�H��ZA��ת�adzr�m'�ޮ����y���_>3qyV��8�w��%;@��e3mE�4f�|��(t�`��=:���\�=���A�}���������Ի��:��=�F�3{)�CE.h��/�J{�|EsW<�bE��$I�U����$��W�H��*�V���~K*���Ð�D�N=<���,Y����=�}>?d#�j74����2oĳ	���xP>�@�D�5^�c(����;���8�cH<�x{��6��Y��#b��O��6s��I�.�	�;/��A�(�/fPg�ZƎ_����/���u�Uc���Nx��ɬ�C��wn�k=�-������fI��p�؊�]���"��:-GS��C���$2OL�:)����r4L��� ��?If�Ҥ�o�0�=ƹ� ��5$N3U;j�),����P�
�;���u�n��+�AG0U
I�abڶ"K��f\#*@����C��B�k]�%<�Gc~q����9��4@-#)B��d�����L����U����\����گ���?mL�Z_f󂨺��H�O�wa��v�ٱ�Y���壁�����m��$VZI�91�cٸ�Ηvq{x�X1�{��%�K�´>Tl^�)ޠz�*1ϵk��4̲XlxVHYEB    4b7d    1310cE� D�	�I��ty�A�+��;�9TQ�u���1��K�7H�G��&�\@N0��}1RJ���C�j��xko��c�C]�m�n�t��KUG6��-�~c���ɡo�����-���y�����s�V��=�4��M�h!���p:�&3�����w��fA7���O�q"�o���}>�"�<!p$qk��/��z�Rn��E�[.�⁇Nh��f�;m���81)�`z��Y.̇$J��2M�z{\��Q� ��Y	cɖ�HI�J�=�����G(Jx1#�䚄�3ł�z���$K��L���>�z�IH2%��p��X�-?wL�)� L�d�C"J��HJy����Ί8���t|M@I��t����R���z� |�-݈�/���=2�K �)�\)d$;�F.Mw��+�#��j��VN�����_l�!��䖴'�7#ɸ�;�vE�[�D�ۄ���B[N�$M�Rβ�o�QRt(�)���h���p�5%��;N�~�ė�,�g�&e{L!�����(�;�a��XK�AG�eu(:4�Dęw�_g���w�!��%�ݬ���-�� B�����P�ưݸ7�H����ဗ�c�؎��O�"bsa=}�q�  ��bHn���/�ֈ��J�^Vp���M�	)Q3���&#���g��I��]�<ǘ��~�T�����gF.��R��?a4p�A �f~��TW�~`�m9c���%94�q��!~�di]�]�/,�Q�0��~���
����R̫�_t�W�\
����i,�
HqW��,����4��'w���)c���y@���8=�T�SݿY�'5�Jc=%�01ς�
Z�����s+8 ���iFc��q��,�����u�}#�w�.���uR�sN36F �5���J:���mJ��et��v��:XTN�v��*����P��%r���V����5m�κ���o*�r��\�8*��qY�q�2�k�6�f������O�/���p�`ruX-���4ݳ�%R1���\�+^�����mz,M�B��:q�/���D~2��������-��z��F�أS_ud����7�I�Iĩˁ�Y��Ȇa�
Y���`�'8��V�<qc�wFoYn���m;��@�rvh��V�C=^ݾ�K�l_�d87�}�ర"^#���%��Jq�#rM_�7��k�<zY�7�JjUr�t5��ӧ��?<R�(5&��ǂ2z1��+w���3,��I�y�;+Wq�c1'�:��{����\����Ml
�J�+�m��a�
e�1c��@f�l�j*�gR0�le�xW3�>ƣ�z�w/�Gd`+���\(�U��&wo~�hF���!	���Q��:�\��⃀��y�#!.}	���`bu�Ӓ��
snY�H�]L�W��p�7ⱷɁ�TL�.��B0�tYwhp �P�����&0֛;�1m�����@-2P�se�X��1�7�6�`ܓ��:�-f-2a��αh����sJ��]�f��������荟�:�)�����&8{�Q����J�rw�*��!�68Rb��T��<P7I�α�Ɯ4\T�-��s�m�(��ɹ]�%&�!O��A��W9o�-Ms��ӗl�:��V��]��i�O�����@5��Bʴ3�u�]�?#d1�Dֽ�_��n�W<D��oG�t��(���)k��*yfXɲ�F��uHq?݆��� �FPoHm�ΗƫEm��9+�&��ǑY��"�=��g��s�w�hZ�lR�5P���+�W�C�9;+���8XM����S����x)�n�
w���.c�|p,YXF]A+�%�?�\(��7��_8>y_�y�QJ_��t����=M>���H�C�D3�������W8�#��C�̠� ������zv^��5� �}�M��~�L�����(���I�X�9�'R�l�b�&�}u��%��kq�����΍�0�A�(��݌�!���|__��,V�PB\Q���J��I����v��c�ٖv�dd��6�u���"�d����.:�ʅ�������I[gr���(X������� ���\�bh�6T�V%P�0:�(�Z�V
I�{;���(¥�GI:2fZ%�D߿vP�X���TT�s��L؎N��Au�!��?C�;ʃ��	7L
P3ϟ��}v���l�%	��Lo�R=��B8>�<��E���bA��䵕U4�_!*�#2���_`�z�����M=��F��OZ�A]F�p��4�����I��I}`w��Fv\�������eLa�)�WL��w���(x4�&(p�b��\vȣ��ք�Pݫ�{���uNe^�h=��o
B�o���K0�4�7+,놥:z��p�Pk���sFp��`S��
A����%{��ga�����_����˻���ԈB�%��j�D�R(�d�b e
gJQ�n�!Ӄ�p��m��x0$Ou6��s����F}��O��a`���O�`�_�H�f�;ԘN+���?x�E$i$[s��>[��c_�
��d��J����[�|ml,��g��
V=�����=��� }�@�-0(E�Sl|�nt�IwOl:t�#tB���Fb��M��	��V�U�d�cծ�޺E�U�y�����*=88�5a��xmG����(i�ͳ3ulL���G.�,D�U`ݱA�E��ae��e�	_
Ǜ*��cJ�5�e��_���I��.s������н7QB-�o�:&�����|��Rv4�x��xj,���s˵��r�D~���������`Y�������Ő�K|�ē�--F��z�A24�XN;�G�]1>���K�m\�h��W;v�ڲX~z�K�2�B�R�W�-5�MleLv,q��h��C�C����'|	O�1u���Љ�tI��e�1�A\E����nHqӽ�eCh�{@�gs� �ȉ�D5�I�@�W������1<��4tx�r�k
����η��7�S����������A��āg̃vl�/s�C��[xc�f<fTlҢ�ao�����h+�l���Y�9���t�Y��I(�����[��G��kD
�lȌGqp���R�+4¢��t2?8�jܝ2ʚZ�0F�X1	9�A�ZJB�M��k���M��.s�<䉐SX��]?:��k����\/N�Ue�©�%�m�!��8z<P�_�=�m��QO[#�e�"h��fٖ�X4�(��@0c��t�3�5�9�[;	�@�?�sxz���.U�2�&�m�yeNU%Q_ܙ�������(#�ưe�ٯ��~�U��=W���5�T�i�2�j'�� DZ�$I�~p� 詵���U��X���"sL�|�/p���F�A�Mኯx����f�ۢ��mQ�L��<���a���O:���Y,�Ќ����}��y0OV�����sQJOg���ٸǽ�=��c{���EI�9؍���44��kv�S��"�3�b뗑^���v冷�;��
t�V�v�H���@�I̔o�D��c׿�d����ӱ���-�t1*���	��@	�� Pt'=F�5J��P{sG�mj��q�c���b���˝��aY�����IX�����8� 4N,d��A�����=AR�,��2���z����N��Nr'����*$5)��������.�)��#4=���A.��id�q�
�:��!�����"�)�2���;���1E� ��'F��V��K��:R���� �R)��`�x׈ ��Ė2�S��qⶭyY-ret:X@�'}�N���ö&�y"�x����:�z �<\���U��KZ���$�P�8fϸ�|��z�]��T,�#�w����f+���J-�Fן=Ih�~���(�w)oW�&c(����%{a�V~`�k�87)��K���K]Mo$*`z�Σ��6��I~� 7��I�diυ4�dI�
BN��5�]'bk�ɷ�6j��SINz���
���ٲ.rZߧZe���2��� �`�$ِ8�9"��F��(E�x;�ӞeDL	G��u���@v���UZ�O��
m��T�V��\��e $�دx����`G[��8&W%�
�_��c{(��B)���s��q `�3��7�S�=�Y�X9J����C���|X����&�^}���S;����Ʉ�h���N�/����7&P����+.DڎQ��K�eC>1�`1������)LŒ�@��xUtك`i�oM!
�� Ƽx،,h�H�O�W�F.�:�d���&�p��f-�s�.�89�� �c�~���k��c$��I�B~�Pt����T���=q�r�v��0����T��7�c��y/p-4��0_�D��ZWSl������ˠ����\U�^¬+��Gڜ�o�S��ׂ��!ݨ�&���dLj�P�!A�䏪6�Zr����,����T�*�}��^� ��'�Nl��e*'�	OXq�ݏ��9� �F���Rx}���B\�­�\�6J�.�J�B��o�[���1��Bp�G�6)-|=���M�t�e�mHwzs�;���&+���}��-a�K
�'zJ�-rH�q�1Қ�ӕ�%�)��1e���u�'f��~� \��P����p��(�Gi��XY�y�	�a��Dı��Z��iE$�A��7�#Q�i�߻2���[A�G:����^ ±�Kn��R������jn�H�k"ތZ�hח{�8@Yu
�D�{��E�7����FZez�� �8��^���3vW�;/�*<��Ӿ��5�sʌ�f�>Q.��������