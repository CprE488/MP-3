XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���t8a5&i?�+#�׼������H���eL*${��w ��O���ȝ9�(��Wm�x���9n��*��)1���>��s���4���;�*y�K���,ĕ9�.>\�d�4U�2FX��y@�*?��@}����1� <���>l��M�܋����D�T:��Q���n��(�Ǽ"<�L��H4(NH�/YRF$�5ܨJ�6�fE5ig*�����'���M�Gg��NQ$�W�SdC�+#1�<_.u�����KQ��=�qe��%�e��(F��B�Uh�.�V�ҷ�Z�'lGM���|����MV�,�\Ō~l�ނg�G޳G� ߝ��~���ϞyH[����.bX�v�AԬ߻�\��.2��&�����L��L��V�S�y��>�\�J=���ɳn�|�kr�#�1ĭ��ǈ���1*I�K��'���F�T���R��ߡ���҉eJ�l�AM�~2*}8a	$\�L�ױ��a#��;�^�Z����2�����7;��	tRi�we,�[F��f�Aaaf (�7Uk�|s��{�@�M�E��f5Z���ٹ�����-GG�����$i5�Y?��ss8W$�B�SryK�	���P2�L��*R������w&1�4M�yO@��#M��a�%�5�hf񴧙y�Iv�1I�5�:4�Md����T~��<���"�¹�m�+�n�	C�,���0�p���d%)V�"��Q"��0����D��`�m�����:|1��)�iF�$�x�l|�)DXlxVHYEB    374e     ea0ߜ���:O�uFR�r����:�e9������[�!�Lܞ� ��~�M�%����z	�h��N^&�+A�rBѵ7|9�E�q�iR-�p�>۲��m6J�-INC��u<2���5�-�՜��N)�u"[�d���CН�+p�]a4k �Q~ ���2��+�ۅ@�P�Գ�@���6͜�	��+y2��'������]�f�:���6�0��S�L$Wt�۽(�KVʖQu	t��LQv�J5�b���I��ܑ����($�yR^��G~t�w_K L���Ǜ�l/�C7D9����!�,�+���j�<��+�A®�q�Ԉ����tA���찍:`xJ�ч<k�T���+��:��'A�J.�d ��P#Vɚcml�ʒd�`�z��|o6���J�:6j��A{M����RUƁ��@;�;��k�⥇/Y���9tڡ���ɱ�!���+����C�ץ����
[v��{�L^�z��oi.)a�([Ԣ�d���M1��g4\0v��J������=�&�Y�BO	�� �TZ��]����c�����l�O��q�i�!d0��O�	aW�\=5.�Xi"�������"�!󑳪�v�T4��KQ{���?h��N�������u��p@bk'�v�":�=u�k��r�n�C�ܾ���yr�zR��Y�Z���A��w0'�P	�C!���߅<�{���}�-$$+�W���)�B5��:�hy*��M�>�P�7�L��y��z��q/�Ǳ�g��:�)I.�U���2���������u���s|�x�ϯu�E�z��ei�Hc/܅��,��n�(7�P����r��8�D�*���Z�¶���iC%�T�0�-�x�˘lv�p����@;��EA�;{R���w��s̛�i�]|�EsL1���X��]�~�:�f�Z���GW y��֧�^��j�_}��EEM��@+6����N�Dd�V+'�k�==zg�Y�Ӡ?[���g�Z���`�s����?�{��w.�H��Bi�P+{F��J5��H '�H'"X](�,`���%��C!`C��\�1s����v*�I�t�!�=a�� �ҟq�����������wWI�C.���q-Z������3��.�����0���ĵ�%���K^Z^wd�r�rRy��>g8��=�@���7>F>ɯ�1�֢��u�����fx�Z(�R�t,P�k�i�_늇���u�~���e���!k�'5��C�������5'̛�7j,̊�R����d�dl�����狑��]��=�DG�p�-����紳�~h`d����1����k����0E6��K�x}�Zp8���<������?1+)a>�|�U�6�Y	���3�j�
�2�#2��oT�t~������5��?~�~��G�}�^AS��A�ڝo|��������fg� ?G�
�����y��1L��T?�yv|:�M�"6�K�#c��٠G�D1���$��j�x�S���R|(=����	' �x#�?���3.۶�Iz9rԛ���ށtZ��e���d,ʏ�b�g��n��x(5�}[:��Ϸ�N*�-�������m�ayg'�JWgN��gd�թ������0�(ؼ�g���<�>v]S78�{�s�)�*��2&��C���(���^����p�~�V(��2��ת��춮���� ?�S@���)x6�'�傯5=~�/t�y)�6�����#͌L6���H�Q�2�����M� �,K��:S�{ck�$ܢ��rS�l�F*�
�>&+zY�\6L:�.?����҂r��AR�oh%�W��&E��'��������eX38K�Y
�׬�b��Gf���ь��p�$4�+��\�5n�F핢�_�%	m�>���Ǆ�������E;��%_��lm�Q�D�Ԭ�M���Rm"c���&r�k�췊�uE5o��@_m2���q����4�Q�dH��������=�K-�~�5�! 2
(>�
���d�}}�c�E#�i�X�>�̙�Q�RR����{ ��E�1r2�C8%$j��o'U5{CP�}ث��)�Qz�Je,L�j�u�t� A�$�gUQ,��H��v\9��I�!R۶��)k�����r���˦��c�M�@QMȾ5���r�J�o����r��H�D9ɳ���U|F�8E�ax_t7	s)!z4)�%Kj�.��g�,.V��0�3���ZH�0�h(ڍg�����Jm~���n�.ҶH���	�l;1a���2-w�)�	*�'�O�;9�%�7��p7)�p�a/"�	��0Ru/�j�S����b���"\G�n���iʵ	!�Cn$,P�{���H�ح��.(�;�J8t�y�Qu��G9[��8�e8�i�r<��4z�1Ӛ�8E�q ;����J� _�o�6����/��&$�J�g�b���|`���ǅL��#���m��U�bQ�yI����
Vq�y��n?���7���Q7$lD��Fo��'�N���"�C�hKpZsv�5�4vf����$�E*���O����o~��'��C�I�P�H�е1Ϸ�#-��Ft1�n�/�F4m}�_�''�vK�Ьx�W�<4 Ӥ�b'{8YD�}&�Ӟw����hD��X��h?�I�l�x��{���EW�%��pэ��6x�8ۀ�B��P�,(iӁKm�ff�����z��q,�O���p9/P�C��L�SS�̊:y�~�u����uA�
v����g����9��.Eh�SY54�zX�"��j�uh֟K��;����	����� q/���2).	ns/�
G8D�,�`V�*ZhŢ�(/��7�=����'��p���{�;ҀP���E�Y�D<�t�(������3���+k����F�c~#��O�� r��b��p�%�z#�D���^�,:1��s�!4
��k�xz���i��b��c��%�>����H����cb�������j��ˊ���4��ƒ�\����@���kB��Vk ��+�a���$�b4���H ��Z~J6��f	P�u4
 M-kd�ID����9�O<zoV�@�����'a���d�ش�r�"�	�qp�^i;}G��?H��P2�}l,��B
tT�ѨN0��ϡ��ԁ��*ǵ��D*�̊DM�1���:��(W^/a������		v����B>�Z�o��������M35���։������޻��0�q!��L-J��v�����M�-�����/��g%�i$/FH,��#�B�Dkg��k�L��d{޿f� 6�	�X�퀾!�k^�7�m�6��� r�n�q7��ѵ�Gt����FO�����Z����iH�m���`2��p��q��u�r�y\n�7��B=U@U��BN��j�)Ў�_������\H���0++AH2���I�� ��#8S�R���=�4p���G���
���X�`OH]�.W�%��L�b�kF�hȒNv��o�on\�!�BM�`c򵊦�j�q�aF���J�2�j@c��Y�LS4A��-�L�S�ߊJ�8^[�H�%�s�`�F霰B]�����4�5��pA�)ճWX������¨M.ua�_e2�����i�_��f~{iD�g�b"�eT�W��܂��>��dM�	�W�ľ1^,