XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���������l��?6lM�q�����1����Ļ���a� �M���=��5ܮx\�G���F�Hh���:d�밞w��Ù�NmR-I�܆W'�_�BMrQ����\� NQ�0���v2p��x�\�d<�ĭ�=�,��*��]�_���S �������G&	��O_*��[{�RE�<�7z�s��o��8�D�	�s��Bv��v����H�=Dˢ���8����A�/M�7"OX�Ҳ�ŇTm�δ�a�����ir��^��]$����8��ٓ:�DN�e��k��	�ti�{���S����:�fbV �3��RBd�����*�y���+��n�g�r��~=e�g]�s
������mh[��;�	�ˀ�@¦2j�#ä����&��J%�`�2�o��1�l>�]T�C�{N�7��s5�>�v�m���4՝G��\�*�#5�=	�Ts#ۿ5I΃�5��"�^6ܟZ���H쀭sa��$H?�<E�x)��3ޏu���2�YEv�
�������V+ku�`h�q�K�2!V+!t�����	��U����	����w��v�����mlox���L��l���IdA�3�������#�h���6���@K��W�W���\�RJ�QM$�6���v�|865~Ll�)�״=Z�����)a��7� ��C�e��'�e�8��C�l՞ꔧ�����UL�����v Q��b���'Z��MK�{����q��XlxVHYEB    7265    1660�*g@ksDLS5�뽳�_9:�(A:x��}W�Y	%]�1�n��Vb�k��@0���̵����7���|U�@F��[#��9u3��Q�i�5mm��N��l�\Nh� ���n��!c�L�.��.���/A���p3�yT�.|#]�Ҙ�*�u��m�y|�%�g%�W��fPd�}�S^�~��u�D���J�����J�^3GN�a�Dɷ��%����=r�`�ܥ�V�mR�3����#�h=�����W���]�s��`��յW\�h��l����HN��+���O^a5��\8��� VN5�t��ZO}8~B��{>�Gk�7���/xi�&��A�=�Jڳ|HTa�{��WB�� �#[�I�;�IE��'�Gy'��ܕ)���UO�@�#ej#O��z�e�HL2:-ς��_.�X���?z�(8�K��cE�<f�����r�+��t�Ɩ�"�}>9b�^�uDcۗkg��չla�U����O����zNx����f�L��1�`Gñ�q���"	%⨫�UK�WcUޔ��"(;K�΁�?�e�G��v�W�%m0�t��"��r¶<%u[z4s��D49��K�����i��"��BA��X��9�EP��F9nݥ�|�L>�E��5�s�k䎝��e���'uIi�h~M�0A�ƚ�2�=0ӷL�C0�d�O ���ř&)�Ge_��,����PC�$G	H��H�:|�G�ur��g>/Y6�aoe�	���/�s� ��
�_Lc�:[/�0I���"�<�<��=v�ט�Fr���Oϑތw�A��>n�d �p����9"�����h�G���j4,]�t�Lq6B�r�UO_(r�Υ� ����<�"|��Eo8��+߂��GAZ|��@�ˡ�tu��G��i���C:ġ����?7z��D_��b��(D8A���d]�3���<�� 0��ׯč"�_�K4e�m���"P
���Q~��ʥo��p��4�2�B��,�%Q�p�V�aE�=tk�?���������u�G]�3��S�*�J.{��L�5��3���ѣZ}6v#��ׯ\�&)�{��:�ų[DM����V�]��T̉����s@��
��dԲ��;3;���a1'���Xy�������4�d-��a)B�ET�7�c�d	I��G;�D#L#`㼎��a6�O��-���΄���_�	��{з�?����&�?�?A��u�՘�p�s���=4冄�Ԥ�?]�N���ݽwR��6�nrm�гJu��<���ٗ�ω}��U1
��-�.T'��-�y0���MzIe\9��!d�/%�.�u'ٗhr�I�����7�cv�z�k��1��� ���9���I໏
!�&	8�=?��+@��^���Z͚�h�l�.h�����\�z:u{tMSd����>֧���2�<v�q�B�ɤ.�H.��(cR<q_ϘU��]VI��*�i�t�0H;��R�嫶����;�sy��0<}��(���n�)��d�L����Lr{b�m[0^�SI3"ۇ��x��Rn�q�L-����Q��4B�<��:5��OO�[�a\�,Q55����W�`=>����O�<���3�*S���S6o*l�_v��QvPE��*��F�m��3�&��e4cK�ױD��7b'j׉��ł�x�.yl�r���8�bBῷ�����9��#���J��ަP�����t=���;�s�܂)�`f��n����2��B
����6%q�R%�%�=�:�E�P��5h�jj�T]ϝ��CP(�O~7Yyy�������q�(�I%/kg��PM�1�WƵ����s"�֕�<T�yyA�}M+ޏ���m��65[~��+]������0e�����3�U��a�iJ��m�!LxTku�{V&�k����{��@qWX$ZR���q�=��!�اQ(�&L�pC�!�ҶȜ��N�ܚfnJJ̎xs�-���1�-�˥hUH�?�Ƀy6��GA:���u�����z^�|�sKN$y	1<��X�ԉg,ei��A�h^]��H�σ��m�/�xnǼؾ�{$N�O����`���9���U������W��(����Y6�A!���'f+jz�Q}PَX?)
�T�F��JT7��dTl�Fdה��%Uj=�e%��;w�NbH�jCჶ�0}�A����Z#~��%d1}��!��j%z�黝f�����'~+�~��g���<vVݯ��K6>�b�+�Kz%�0��N���D3����\^�M�OÚx�po�1�1e�$���4y��)ϙ�w�Q��wm�fU�����E�O�t����Q��.Ѧ��J��CבFl���̢�WMT(�1b	YcS�2ں�/yV����;�+�3�L^��5E�*2�!�Ś�-ncV]������	*n�{�@�����+>od�ڜV�<X��Ƌ�R�������o�C=-���gq �C�t	������/<��%�8e���=b�Sӻ!U4e�0>��z��"�rct�8�W~UHK>Ƭn`s��,4�Y�ث�G�q���@����<�V(���թ*�];g��,�GEe�F4��!8e�ŭ!�z�m��k��!���ギ��X��?08�[m�aC��\�'$	��?���޳
�8pI��<�=���=ԋo���5e���1r4#&x&�w�����z�Z
'����?�%�X`�k.#�B?��TR3���5�PXz� �x(�Y�|e������.X퍽���P
T}�c�Ï������4[���Ǧ�Y�2���d�P\*|-|���EcֈX�8�t�o�d����4DI���C��w)��#Y
��BJ8������ R<2�,>��0�0������,-�%����O�����m�r�6����8?��E���%op�C�ǲc����i~Y|���R�v�y(P٣<��Nֿ��Q��ܓ���F&�Z�\��ډ0��RR�Z���O�������8��_pl��mh�,��	�Vc��w����^Y���d�⇡�ep`�����[a�brq�Ьl���DH���8���z��;��s�E}��E5�U�WhDܠ�S9$"�F?/�w<Ȁ�����g�8	�Yz?��(�@�SWm%�L9����2�"�*^�G<\Τ9
���Pj��V���ʠ]l�%#����"Ⱥ�'������h�2*^/�l��ߒ5=��Uyݫl8)f�ں��EL��
g�1l��5
�IN,��]�m�x[���
ktʺ�F��M~�d
���+D�S���A('2�b���̵�+@� ��~�N|w}i��t���1��uwe�(�f�(2�����a)'0�!~�>���R����ɳ����6L�$-��1�����Ҙ`w�X�N�� )�hi�W��gn�:��c9�5�` �+��$M���zf7��+"V��jn4>j�e����-���<X��q�'�K߉6[5j8H=�?��i^����?*0�2��0�B8r=�xn���%�yʃ�����)�f���#t��:)�F�O�r��x�����g�ur���X�{��\"���T����-�x������'�z�� U�9 M�F�l�z&ٻ�0Tr�*:��Ə)�W�����4�ZN�E�Y+��A�y���ً�JwIB�����A%j�2C_|��97��s�`k<�l�Ta��fa�C&j�`����nŉͦ�W�a�D�3z�&\�DF�i����
�9<:Nr{�	���0���!@�Cr��r���S9�
[V����?6n�ji��]h8l�����T�"���2��:���,M䈋ᜮG��w\dْz����!Y�am�0�0d�\��(j�ͺy"�kCH�1��Kثz�ӡ���r�n�J�� 5�����3v;`��Պ�sf���
�B�
�ҏ��Q���d|�����
�7�nͳ�!."�)�*���.��d9�&EYb�1Á��]��ж�8b�m�h�2Fl%J�����X��9Hx�֦��n�	�@Px�y���02Uh�������b����H	/�%�d�yh����?��0��g��Y��g���y2H�Q?����umzRh�y���=Jj�2��am��M:ή��_�{��C��:^c:�|�p=x���(SׄK�H�q�qp��JB�͖<c�E�=�����x[�]tqS�ڭ:�9���N(��k��.�	�C����a0S@Г�9�ɫ�� ��Kq?�������e�ۍ�ą��$�?�x�:7`O���)n!�?��2�� �i e�s�f xv(��ÊU��󚝓SA"�a� T�#���N��ë�i>��W��@9�Kb�?���2	�e�5W�cSi���鼅w����\Q���.�7hs���(f��Kv+����:D}�ε^�+�i����M�#���a��4�O�2�:D�^�����l��7�	�������3?�]ݚu�� ��Kv����s.<��m����1�U���ᗜ9��udҹ4�� /�Ѭ�{����^h6z1^��F�{mU�
�'��4��(	 "�|!���2HHBF�$A���[��ԫ���Z��x��;��0.�®���1xw���`��&�f��H� G
O��tƍp', KI��[1��K���	k	����BO*��D��S?�>8�X��Ħ<�F@_�|�_�Ϣ�L��:µ�v�fĹ�ѤM�JV�H�ޗ�hs���o��w��r�kl���p��ֆ�o��?��s8�1�i�\�7:���F�i�װsh�������\E�)���N!�0��KvI�m?aGf(a�X8��\�t�^�T$���id�9_��d7���ܩ���ߕ�X����7�X[�Z?�%�m����Q΋�Pئ�Ӟ5�Aoz��ȕ�y5SBba�>�G��O�`������莻>�	���mF٩GΪ�Į�/���$�����i�ٱ�$��=�?�#�r�k1<���. �{;�	ÝU�2�R�5tW�J���r�[�+ň��Q>Sx�<�&�HV����`j�V����U��'����nF���:0�rZ-���U�&_q�]�Xm;/g�A9�䫤7>��ӌd\7�@v�������4r2�).�=�t_���# �GglT���!X��bL�oZ}f�8@���Z�0����(du��2�"�7��p)�A���aX�p�Jˏ���8�������r��οǻ���z�*�����W�
����7c�@��hu6���:�1���gd"C�k"��U.2}G9XI�PA�E�?n\���e�♲]ŚJ�T&���8��̞ȗ�!S�՞hM�2
�}SÄXq&����Hp�&�yd?bߖ��ѱ�����8��
dB��c���]��ټ9��L��L^��~'=�,�x��0vy�%Vr)=�R��]e>L�Ð�PFUۼ�0�����_���7ˌ��~W��@�%O@��DR4Or5�+b(c��*�J�N��i<D�'�^mk�9[��D�BY7�%^Z�����ok�/���rI��|c�r'�+�	��!�̥31�(�t˲@��6