XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������/�5b7l[#��M�8C�^���}�u�E5�g<��qBgN�9����F�O�p��	��ơ�,ȶ��O�YM�Q���*hC��x�y���ѝ���"N�P�_k�lǗICW:�*�@:�еbԃ%��2����<�G��=����D*'����k�'��W;� "�L�U�.�����8�_)C�����pr���J���r.{��q��Ȗ�/s1��h����
wp�+��k�z��?���']��\�L ��#��fr�ʢ�-{f'رO�S벐g��p`W�o�6$ki=�8p�ha�+?�8�I;��W�-ʳNR�a���/�,fA�YM� v�cdC���)}u�؆��: ^q��C�� �C�������U���S�s����egQ�@�w�}8C�#H�ThuN�o�-�`��8�2q��gĔw{�\JY��MW[S�E�ܹ?l��uS��"���}�N~�lS�;%/�O�i'֎4�aZ
�#K�c�)�J���<|�^�Mz`zz{Ҥ5-%��?�g���������{�<��>�9X�Nm�*1���oR�o�ٖ�F6v	e�6���便��v���#�6#S�������t8Q~(x�h ��Eämz5��f�[�j��b������:y�ZY�=^yI���|bLƸ *�*Cb���j���~3o�d��0��8\U�Nn��հ/IQi��L�sry\�=�tE��-��� G�?��]�dO�:Y���=i|�Ί@�g@��]4��XlxVHYEB    4052    10f0�;Xd��nrЧ��䧻���$�/��-���"����������K�8���E]�:�]�]�yP�肨C�I��Ǜ�$Ѯ9�ۮo�M���ZX���~*h�*\�j@��g�^jH�}�S��*��2)&���>J�G�� �8���-\�Y� j�P�������`�@r����	�h��f0Tq>���?+)1y3��Z�̓��n��r�6�ISe/|-"� �}D#�~�/ƕʖ����c���8�;��"�̩Ug��k:�k&����g�[��ՠ(�ޙ���+Ȧ�(6�K�1(~�8��ޱ�ڧL���%�9�����%i�'��!kz/!���� ������pD-2�2��3��{�u��ܢ��EUh'�8�x)��Ѝ
4;i:*���^-�L �UerEw����M��+�zש�S81��,���~v��q�XK)��V�ƇvV��dW�̥��v��ީ��OD6.�6�;U�Ubs\M"�>��op�җ�!7�t�r����k����h����)@�fL8��in9���p,�R�����k[K���cùN�H��t|�:�)0F1>�@���j�/@��
�c�~9D��7<������� �3#��_,�ð����@pn��1ee�x��}D��n�=������jRqT�1��N��&Üʅ'���zhe��6�x�i`�l`˸o�>��cfr�F3�)���4����F#��a�8�3ެ�*1��j{d�Hg��v%��tnqh�iL�� &p��,�*�4�:|S�@#�P"�ȓl��6�\���Br�lm�:��-+����JO�)4�uN���_�Y�bb7�Eʃ.�]
=o#��;�BQ�`���{T���U\h���T?�u�.ԡG�$+�;�4V�ЭC���}�e[c��ӄ���y�13��Yƒ�f�ͪ��q��4��s|����ih�������w;���B�v�7�,g︡ M0JL�s��[=�>X�f��+��RD�q4y�[���bo�1!��Q6�$F�>�Ɖ'p��6`��~� ~0��&��B۸�H��qY�C"�M�F�6)�a�ԅ8R��<�7Je(Z5�4��Bx�n��2�qu�K��3��jDt��0U»��7�{e�����.K6���~�o�o�L����P:^�3�`�W9�������U������+	Qekl��	���*5�O�������/�r��E��>pk
̤��yWeB'5��06��<*ؾ1[�m�M�d@ZD����Y�;�Tw��b*|�Q���E�%n�	��`�k�����׫��,؁�=ʔu�jš�6�O�9CH��^��k,��G�X�~2N $�R�������&�D�P`�M�
կҿKQ�]j'�y�7��sT�gp
�
��̓��<H�B63�0���>�P�wr�cöxF(�E]���V�VzΓ[�fS�L;�t٥�Cz������(��!�u�9ɂ�N�	I y:Ҳ�r��vq��odc�V�1��m��/���G��W;�| �� �z��~OB?Ȅ���B1'ũF��$
�gt�T��j�	4����z���&�����e`#�mG�k��i�AGb�7���ۼ\�?�c�χy]X<��L�7,/Qg�`<'8�|m�|5�[S6>��ΰ\�-V�>)W��Z�L�lW�K��r�%M�R�4;ܙ�1,r�8׶iѲ��!�t;�dw�d�}Y�K5M��R������������=��WH]�H�3��w�jw�F��?:��xD�¶DS�7�dv�S<��P����LЅ����?�]�)��A�;\6�ז-d�R�@�nl�+�2=�YΤ����mY�	,3���a���ˊ���s.�y�Y`O�`nST� �(.�szq�'��TFU�Cx���z�է<�׋u��V��!�2���[��@DM,��-B�v
i��Dl1h�P�[>x�N�<󑗁H�&���4�%�G9~8�aߣ�OO��f��cQV�w�HN�]IujÀ�굖��E���ǈl�+�b8B0(�\�˒*0"����߬X��@�q��fT���툯gИ��EB����pb�V�ͺ|�+r�lµӲ#�y۶n�Tb�9K)�I{�|�%��0E���C����o���������G�7�V~��lVN�D6���vK>�Y@Ӎ�*�q���20�2e�yG���̤�������;;w$�˶(�_��J�Ԓ{���wH�0�4'�^{7�޲�dkwm�;2�?	�Q_]�Y)qOK��K0H'��B�bN�=v�� �?���<�sGٜ)��s�r�?ִ���w�!���/��A'2mIf����-r��\,UfE3��tK7�]�0�����u�:�#bO��Ʋ��-��yPDa-��\��NA�[�v_��ϋ_!��W�
�k}�E����Q���mx]�� w�`����tu���\_���_��qW)A�a���=<DZi���O�[7����[D�d��ݺJE��U��oa΢_�x�Leщ��P�"� {������ƨ7>��c"8%)����0n��@��)�h���������.9'Y�OxeB	Y5���j�$ўp-�O@��M4���@T����v����T[�nxC������]�K�۳�]�*vtFj���|���M�U|�� ��"by��bNgY!�VrƋ��`U����]t*`�w��t���-��'HK�7��T��^�7n�v�I�42��PXw���3ٿ�n��#$�ݡ�cg�H݉�����M�`Q�������<�"֣^�{�9�P���J�½k�|��jgД��lp�n� �f�_b<�%����ڌ̗4O��^����N�J��*Yb,�X
��� p`,�4V�P�^<^��z'k�ZUi'
��Vh��08fE��+h��	����23ͺ�ʛ[n	]!&[&rC�O|.^�4)q��>>x;#,fF���4�/h2���Ue�r^�%��q�%b���Χ?#��ڹ��PH���Q,�R���/G�F�n諏Vo� ׄ:�20�r�j�s��>0H����܌�	Ceq,v!;k�,�<��/�z��+Al|��3���c���W�t-�p\�h��k��gl[�/��
J���=��6�/E�pe�9d�7��NL-z��y@�lè���v4�V���/Z\�y� 7�՛5��Ub��j��&Y��H;�}H��m�w��["�0�5�!�$7�g��^����]1���Ny�5+��}PxR�I���P���^�\O.�G�?5}]k,��V�q�(�׽��B�6�C]�	��;�GM��C\n[%��=�B�ơ����!V�8e���M���{36uy�Dˉ9 ����fۘ1<+�����-�kl��7^��YX%���$��;W�_�#�E�nͦ�3C�O`:nW#�$���j�$�FW�'��?29\��e�V�o�d!3
X؃IF�d��$ʁ�C�BKc�m.����b��|3�k������ ��1���V�5>2���&�J]�ޯ�/��m������#\��;�T�d9��D�:��)���l�|�I����*0�&���r3�Dk���]�y�T�V�Ɔ�^���>����h; �q��⴮p("a$b5��6N4D��o�"<�n/� 2?7����c�{�2f�à7�o`�Q�����QK}-�*�N�┅��AP��w�4<���������h����;)���Qڍ[{v��ȔM�M��'�z�|S��<�d��R�@����o�T_��+�7ZRѥ��y��Z�T�Ch�q��~Z�ݿ5�D�i4��x��C��u/ĳJ�r&E��'�	��n���%�>CGx��8�'�b0'�	�6�-�"��3D�Q1�;��HD�;�h`|)�����Ǆr�Wmru�į���E�!�/�[U��#┐8h/�X=�|q�~Tm*|f��8��O�Q~�Fj"'+�
��2>o<a�b�ő��'�;�B�<��3�}E�xG��:*�}e�@��	��~�-�u��_6'�N�B���,JT,j�m1�Rd~�����Q�ܫwn��@^�vu����]��@Є���S��V�J�8j�$5��	��:[��"4s�����m�b�H����i���@=�.��@���&)l["�>W�0Άj��[�cX����͛Y� >���A��&���K�Q��{X7�!�/���]�'>��mfΓx��LS��{W'8�Ah=�M