XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��,J,�@�����.�bG��-S��A��7+@?+�+)=����b�� 5%�mߪ�Zgв�rq�sb��􇺔H:��i�?wA*¸jq�;���b0�K߻hU��+5�W�\���?sҝ>ۡ��ԡ%�p��{�V���2q�%��y��[l�����OpB��o�N|H���ɤ%l�F,+��+�
��������C���\ �\E��g>����.pN+b��#�j����]L�;_��*��Y��{�
_]N�r�A�vZ�� 9_z{�B�*�%���M5��h�l��I�G���+#��K�8���}���*ք��<��c	E
���h��*+BמM�ڲ��v�sZ]p��:�D�ZvPg �R	U�t'� �[(����b��!F	�Z� R�w����v -�u%W�<���,zj,��ͅ�u�t	e�@�7p�Ԑ(;E"����b�^�&B% ���n��~j%՟�L��
�u� ,H(kֆ�w��YQڿ�{���qKw�����s�o��q;}��m�j(R��$
����������I�T�zXZ\i�ML���B�����n6A6��¹�I)�M����� j�>��W,�V�C�ÜQ]ʧr�w��r��8vN�*q1Ïo���!#ÖY�����Xi8Ģ����0��ǈ�EM��p=��RO&��I���K��W|�ْ��U���r4ts���(���ܵs�f0Sgi����]qJ�����v�Q�˻�̨�i1XlxVHYEB    374e     ea0�J��f9TS+#��b�����F��>��"=��@B��.h�3D�"�'LV�r*o�ewCj�:�������+_��9���Ï2�wUp\Z�^����}+to����m��+�ܹm�8_K�
���D�l���~�(�vs<�s�LR!�gpcv"�h����!&���)u�`���|.B�hىn��y��5�A��WS~���{h�uiSZ��E{O�u_���b��R�U�]ߢ:F�'3t���zN$��b����(�ֳo�!�}�G��\�z����֢ Kn������� ��ӠyK�=v1_AӐ�DV�_��2������U�8��x]A���?�'��1��~�Rr���>UE�Y��C�ctTZ���%�p�;���c0P���[lm&��l�5�� 0I5���P��W�EZ{��� ��H�q�?��{���Rբ͙���$�*'9iy�R�9d���Tnz�J��!���G^���8X���-iX�8�����lu��6I �U����e��9P6(>�6�,�k8 L�5o~����.�P+e�˛�	^�l���ͭ�_
j}�h��Lc`c�.�|.AF��\�wE�چ���e�V#����R���2w�ew��ܪF�@�Gx���E�R ����|Y�O�5���Q�A���o9V�v��]&�-0{�M�	��;?����M(aH-,�м�����!�����**=�O���%á5WjA�,xQ�Ygx�5��R��2������W�u��S>�C7�K�2�͈3�Rx��s��7�xKɵÃrO�i�V�K��cԺ�|��N�c�=���$m��)��9�?����_���h�>�]x�i���:��yԀ�J���Ώ�lZ�?��UD�]ݴ�}�KM�&a{��E!DHhGZ��h���%��f�f:�ݔ�}-�ߨp�67~��h�#h_���e����OW�#��Q	Q�ϣ	�,�V
���X�&��H"-���<`�~����ߛMv)i� w[QA�X�XT�x����ÓP&��q��ݼ�\������q$�u�ϷC����dǏm����e�W�yJd{�~���g�5i���3�3�,��%NH�p��P7��cQ�V������.�z�n�\c��³�������=���4z,k;pi�1<-<5�u��iP{%�c�޵��#���L%�z�f1/E�!#?�ب�=0����ݏ��K#�opu�up�J�6ȴ0qs%���M�ə�׿��Lk�ې^lQ�w�h�B@
Y�S�0�?=��Gh��^3E�	q�߹U.W��% ~�M��f��<5��m��6Q�}"�G�Е����F��tv����ˡ��`Y�wP_�!�����(�Q�fޞBp���Ŗm.��4�3�!�.����y��nQ�t�x�~��y�tMz1�<�����UF�܉��D��ݜ3����;ږ��*��3��:��3a���"�q��F�_Rʘ5�'w:"�*kFƂ�E�F��8_�Ά7ǐq���;�,L(�#�i��߳���0���n?�c͆�����zt5��c�o�ҟ��&=�:�Nv��u������K�|��P^��/2V�FҔJ~�훋T	��#y%�h�kQK\��2�0,�td�����"�A>O�$��Af!˄�4C�+
�=����w~����=��_�l>��S���^� ��K���%C�G���� ��1�ng"e�E�&Fr�t��ل������r��،\�zʿ�y(f���C�?;m?�w�B��:>jh1�>E� a.Ġ�'�1j<xB�T^���j��G6W�a��*�K� ��ڹl���|��O�~$9��x=Pa��ʡ8w+:q7]#��:4+�Eg)����
�Wj�]�(u�@�շ��'�'V����R�P~N���^@�F{-���D���9xv�thI�!S��Gڿը=4)��ыp���Rs�e ������>�h/�̳d��Vz���`���:�|�"�R=��Lll0S�2�-���	S�����tL��"�����X���;�J^ى~�dx 1�\^��QxJr@#��A6r���2��a=1�7�W&_��He�.B��Vt���5���U��<U�!A]��[��1r(,�Kbސ-�GSn�������nCp,l�vMҀ/���]P֓���4rT�9 ? q"n���죂fP��<�Jo���r�P�}W[#KC:ڃ���sZY�B�MV�Ӗs�2�``�3UΙ�� ���E����
#HTLi�/�f9?h]�:mzb��%�u���LC�< l*Y�����An�o[w!�������a��0���SL��} l���x���R��F�w �p�-�8v�����l��U�J�h2��)�kJB�ㇸU%혐��*��d���T�r��S�j�hb:%�Dɰ����6E��0ޛ��3�4��V>�S��-Mfkza�;(G��>�ܝ+���#�g���jսl��B�m� �y �p]����g��Dw��j�B�K(At7w90�O�	>���"�%B7(���D�]a.�&~ؔU��׼r��٩��&�'�o��8���d�
�53�9:�.Z�g��U�[�1��k������kD��?�>I흯#�Rn�������E��q10��^ġ��y_����Zj[*��~V{D��������!t���
�F�PJ���d�oΚ��4<q~v��tB�S�)��^�}]�C?J_0}E���j���Gi'難LQx�n���e
��%�f�Y���p����-��~��˼e�B~�$��_/�:�X%��i,�]��dOP'!
�tcÚ�B��\�L���3�hګ��	'!L7'���
^�����/��ʂI�٘�Iq����6�L�s"�Ɗ0��ć�7�|;
=�ܴ�G _�^�`�!�t�mh�U���0���o/Y [�I�#6U�6�n�6�wJ�uRٛ0��~��*Fy��q����r�����M��yp+�y�[�b
/NX��f{>
��)T_f�dp�͒�6�n-M�a�F�ÿ8ı�Y3�����f�Lմ�����i�r��D����"׬J��T~>f�����\�ʅ1E�7����s{Gt�x �Z�
2�S�;ZB���bTp?�Z���aN�g��p�M��9�Ɩh��,��h�{I2�P������w}OH��G�N[�V�`{?��>a?:M�=O�}��9�Sk3�w�E`W�r	*�Y�"����%@��Ѝ2RHO�7�u��_ͥ�N*��� =ƨvi�n��|�3|��)�IS.	��	��h���T������0��fm}��P�����N�x������g_��I�l�Us�I;���Hc
���!���a����b��YN
<���ɍ<��i�ޢ�&���ϩgд�5i�_Pd7��M�}�Ât���
C��i{"�s�"Z����v}B?�r,v�.5(�O��cP�H��� �C�nnp
�#��U�mn,jd�$<p�:�T'�:���yJl;��iY*��̼�c\cX�C��K�y������	<�̤DU�v����;��H.�o�9w���s���@�H�i��R,w�l�̀��#�j7�ϭ�E� �9��"B;HХ��\Jp@L���'�]hn�`T��{�&ĵQ�C%��,�I&Y�1��mܖ	�7�c�1�幭�����S�wQϢ6����g��l#ңѱ��3