XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��dP���q��nP�����cs���X���'����d1�_��c���\C�N8�`b HS1�W]�&6��i��#�k�MM\�qR!0�3�ɡ���K8�����b�,��;Y7|-
B�.�~Ωc ��X'��cK���m�@]>b̦�n�;�ڿVxu�����L�*�zy"�H��Pu�X��'��R\�n�v��V�~�?@��_^�j�w�{cf��}���N�E�`y�Q,JTy�,�Iȋ֠��Ҙ��A�s۴�2̍�����G,�7��%gj��{Oss�z4�����e��Oނ�*O�����PbU����&cU��\0���hـ	Ł_�y+v'1�>�U1OH��e���vc��ze�XPx��px����="��s_�z���
�n�!���Gj���r��/6��Hp�;��x�����!�5 ��^w��T�*:�6���ú�ޕ������9�z"=���b�J�W|7��'�����4"Z��+��y�a�����H��bNzj�n���_I���������JD��
r�l�*+��0�/��ѷh�m��!�,Yۂ+�P�tAs�ge�AB�ӴC�4��4��O���7��!�+nf��2���ܿ�/=�J�4hZ���Tҽ����eA�'j������s[x������/x��T���R�3/=:d�����I����4p�	�(�
{{�D���Pª�C�u溞��������,%T�'S�P^z�o[�uN��-��'�XlxVHYEB    76a7    17c05�5Em=���^�2yO_��N���oU��C�7,] ������у\��S,| H8�2O�<����ͬ��o�.b%��dو��8X`0�fra{����B+�,�8MW�ꧨn-p�)@�Y8�ܙ8�~�3YY�H�ȹ����찵��(i�8��i��G��=o�Rf�Dj຺#����ˏ�����V �bע��R���^F��6|m�>����O[�N�H�v�4+��v𻔕RYBz�T7Y�AՈ��_�3V}�!���08G��������� ���6�IK��%B�W�AaȠ� ;�/2��c�:�4�dMU,Tc��O��D`N#_�E����j{�7�P}?���ň��HvR:�IsG\	�#'�&��Z��iPڼ����x�	'��C��B)o:��d<����P�����_�����
�8��|S�E�	`�T&���
�%%o�:PE+Ŭ�����dąkV��G�F��k�/&)��*>i�Hgc���ت�/i$a�1ߒ��a;'�p���	沆�!��6S~��Z��;��D�9тCy��8A�o$$���݉M�j�ո��_�!aLb:"�dP:�M)�A��V^~�Wt�	+�8��_	
���N�/��C����x,3kf9&�`$��ќ���iǯ����w�Y&�X��2�Ә���kw^^Ǚ��3}��h�C��zy+S�>"�3�_)A��*��*E�]V�e|�1�r�[���G&˜��Ǫ��ֻ�*�f����*0�$��_����0=�mAq����n��z��|�EX2�t��դ!k�tM�d���iD�Qa���,�N*�ku����1QU-}���x�-�{�;e�X1P?.k�����v��{�C�*:��G�kUUp�Cc��:@��R�
��~�r����z���oi�S��V�E��$�9i���e�"��Ȫv�qn�I��x�����(�Z�/J�1�B�B�iH�$ׯ�Q{����J4��?#z�A��C���_Y#�M%o��h<8�؅�*�&���u���Y`J.�JwCzyk�Y]Qy*����ym��q�uB �%5�x�m4K�X��� ���������A)&�]m��Ρ�T�j �U���Y�ڨ�ɳ�sxS�T�mDΥ9a�д��3��<�@t�C&���_��w�[�7\Bƅ��	Yl�#��+��KU-�̍��V�b@/���|�nK�wE�U^�,~k_�Ѓ��Ȉ��|�B�d̋�Kd��s�I��� 
���@8
�!)�����+�Eu��V���1	�͍ߜ�	�$�Mr϶E�V��@q�������W�L�2Ȍ8
Da�Z%���{��.�#���	���N��� ���.�,�B0u%�hBfze�81�-�d%gy�mW��� ��z#�z7���hX�#��d����=P-�z�!�[��)��	T�e�w�^��	��＜�s���!���}%��nfR�m<����E�ʏ� E:�&���dܑ_)/���E}�h�e�{���L����L~4�κ9�&��ڎ)2�!���LR9��@0<6���8+��b�˨���A�K��L�C3�4E;ƕouN���{U�>!�;��agk&���� 0o�k?��bL��["�Ӌ�|q���u��g>a���2���Pw�����p����E��d7��{�'!֓��5�l�Q̰��a,��f��y��B�����YV���΋�hP7�ڤ?I���|I�.�F��P�I�B�7�г�;����n������f O��p�71�_�;�3${ՙ�������y�5H�"Q���OYI��ƩJ��p��6�$���wpGv�cB�&'87ϻ<��!��������X�"? �i�eV"��sƜ%��:�ɻd̸���
<F}8��q�����p���X���$��n�Q��i��i�cuȒ.=φ�ub@#�s�Þ>�K��*]d���4�W
��U���e8�y�
���Ɓ�ZxS����1 G}%PP?_�r�B�:�[�ͥ��n)�.���Yr��%�
��pKX����c��f-�2�wN��.�K�����]���"@k|7ʹ���/�1a�'?��'g��XjR?�������Vw@ �c
��k�32Rߺ���W�r,�VW���6�s=�§qõ�Ѧ��[�G��Ĺ=�͖j�GC��*�en�ch�t6p�r-�� S����T�Yl�g�ϼ���L�}����T����^;��vq��z��w�.�7��س��Ϥ��h٥ ��X�m���"q���[<Y��ЦE�8�ݲ�v�7��
a���l��&��3r���#��C{����ߙ!����#�ـf�o�I��P֧$��wg�紆���K�(,-B�f\'�/^���Z(�"����,y�gi��ڛ��W{��v�d��lDbT�>z|�[��d2+BXus��I�Wա����6Bw�߭��� ��������d����Y����B�R{��mi�<'��fcȱ�潧��z�ie1gUS0"-��������q@��(���!�x���FS5ŭ��]��twT��V/zоt\"iZ.r���\.G�����Z���~9���[����r�"�]���䪱tQ�-X�찧�u��TD��\�#1��;����uqZ�=�C�FC�Ո.0��`ӵ�ޔ��Pa��!���FC*�d���=�~�SB�mw-���J4m-������m�Xw�n�<���s�[Zb���j��,�oɩ*�������!�����<����'��z��^��Ӊ�ye�[�x �#���:�s%�%��G�X�{1��<2�=��t�G��!�@QS��7(��,Y:��� �^�n����[a˖w��s;����}3��Z?'"��U;�)H�I�d�ҙbl2&���x��~()"AGo�K�9�oU!h.[&iQ��me/������V3�4a������P�+%F%7v~�Cy�.s�`z��Z�~XfX;�(����4�r�^���l���NY�ѵ�Up�ӴrB}1���eX�9�$x��A߬X�4����<�+m�.�8�Cp�Z=4k���������8��������*��I@�D>��V�� .��҂���^dT����p�E[EE��ɯ���{+��N�Y�t�bL=�P��O;����E&�mZu�	�P�-0ҵDi�>�ٟ�/M瀨M�Q♉�+MͦDb(c�MLb��K�?����x��3S���lY�Z7T�:�z�J奍�"�L*͏��E*K@�_jOwq|~���]��"i�������,b��>?�f"=N�9X��dwG����{�ŭ~i'���;������g	�s�R�\�5YC���9��?׆��3� @d�>��A�����j&�& 4��$|v1�O@ld��
éhYڈK�!�H���e�^�}?<P[Y�;Ql��U���&�����\޽���cܵ2
�F���ސ��g�dfs+��>m}�8���øJ6̎7}�_�d��v���68ͬ낅�iq)Ww�7X�ٻ��7F��u��^���"����&���l[�H��s�UzU���l�e�ӎ���k�I��r��'�s��|9څ8�B-g�u�;^X�S�|���i!���?$�pT(���ijVi?rC*������*��l�&���'@2��X��p�]��֮.ho�%4��*F�mC͒���K��A���ǋQ}��E�9��Լ<t =>�����l$��k.w�t����P�C��F�����<�?��3�l:�ox�D���
�����n�u�P#�I�cÝ��k�l��:���Q����g`�d��b�z϶���>�k:�Mk
�R�F��(;���@�߈�jR~�3u�o��O ���$��z��E��j�_�R�k��<z��s��ɍ��t�ͮ�ڏ�Q��(�)���EB�d;s��8Idf�ZUo����FM
X��	��w�zF|���u�:_"��|��c���;���/��U쪚�H�.�P����M��?n�f������|��Cs��<e��<�o����?v����Mx��8�qJ5�i�L��P�YҮ�� P��Or5�y�Z�%.A�"����i�O{0��� �F��[��o���Y�`��i&arBY�����C	�ST��Z�C(J�y�01�p�t㤎8��0!�mNu�v����HN�c�)��'r�����w�=�"���6����� ����ݰȳ�*im�-��o�P��zgv��J�b��9T\��O�{�����Q��	c�<i�$=�r�h�V�/��b�:�B������Ͱ�m��M����	�<���G���afH_�U�W7��<�ӡW<.���?���_=�|JW���hO(��]q���X�`�b��\$�<�E��rUi`�m6b��k�3;�Y!u��h�W��8���M��
���elu�}�p���jG>tZAȿp��²?�4@,
�W��zg�8n�d���������thy�F�of���
���q�6Ҙ)?���]�E#���wH�/'�&��f�3~�u�c�9 ��sF�-1�b>W�9����^_U����1�/ ��ϭZ2܊�7H�G����J�f�����>�!SkSAmn�z7<����eȹ�񶻏���T9��v����t�xΑ�ű����~%�EI�M�U����^y��F�ޞ݅9�����傃�d�q��K+#'�M4s:�m���#q���xJ�o;����yY���O�F�&��ho�Я��O���]u"�,���o�����K�-E?8׫f�nLZu��9�ToWx}�D�m�����׆�|�Y��6�$N+���	&]T�W���2����[�/���'P���z�!a��r�!����+�1��#���h�Z�A)�S�7k�������$i���8����݈��h�iͬ�𘄾��Z����Ŕ��j��t1���4#��Lx��l`�������y)�5��̝'�x��W&��B:W���Ȅm����n�2�X�`��A2*h. ���ȃ�=�3k/���rlKc�r��"���
\P�;���
��Z×��7GΙ!I�&���z��=��J��jY�*�����-^��<�=k>{��QR�*u�=����蒹�%4�z,H�X����	e &��Q�&��6���:������)���� ���_�Y�|��-��ǯ��>MO�=��!b�Z��g��D���;5�
V#F���\*W��Z��X���M��)��6FiLơlk��I���'�@_���Y������h'�����w�?h�J�Y�D��qT�"�� ��e���+*->K���U���N�c�uU���t|Gz;��<�iP��+��:9~�ю�k��uD��`ڴ�N��}c�h]�qh0/d��f��'՗�f��H)V�L�,��0��3���R	����q��4)��
m�!���Y�����E]���`�W�rS	�i-j���ߦ�$kۡ�,E�r̟fs��7�}�KƐ7P7to�R��"�lP��Q���K'7�Z1|�AQ�����h��!*Js��J m����ԙ�`{�������ix���k���*KX�ŵbJZ���f�C�7�+���ｔy��Ѣ��,����c�M��<Nu"��-�֒�S\s�T\�X~<��έ�R0�T��!�� �������L���ٺ�.��vh�u�ᚱ�6�_rƫg΃���D��<4g��)/��r �����Gm�͈`ݟ�����@�=�>�_i��f6��/�#��n��pO)q�R�tq� ��dP��(�ဦ�e~Z	�Xp-4�p琘b����B�c�6�2�*�n�#�O{,��>F��YE� ���tv�?H 3��K&/ �Y�2��u���V��2V �2*M�����q����1�P�ҩ_}�k�X�e;��G)Zt=:�-�&ӛE����U���k��U�oMb4�}��HQx