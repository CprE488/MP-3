XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���+�t��.Bo���
�pu ��y7�}R��|#�Ht���F���>r��u��2��2,әԥ!���]RFy
C���$�շ���Hn���B��,is���z�?�".k��5�c}��`b/z��Z��(�Э�P�z�y�~"[-Լ Z&#��I��[!0Ե`�y4}I�$������~��F	�N�f��,�T*/�>��I����8b�>#���q��ye��B��b�\�TQ�A��p�q�$�*�p�)���~@������v�qYo7��w�avO6k}���quO^����U�f䷆��� 2G�V5�.FW�QL��͇B��&B��]���r��(i���}fy�U�lW�Z�v�*�E��9������������z?07���?? ���^�.	�;1Z׻� 3�f�.�b.�A�[9����*�RR��
gX�z�zF�.L��rk[(K���*�����q��:��L� L��M[��|dO�#Л(==CK�/1Pˢ�X
�#u�!TѻK��u��=̌��̑'Nt���㎓&x*1�_/�۳��$��g��e�F�0�sg�#n<s�)�R(��VV8~"9IB8��㒎���KFn��3�s��A�Y�n�>kXpw3���{5��[*E6�3i�E�)�:��0��B'Co���;��{�ҲV�n�ו�Vh�A��lc�-b|۪�XL�	Ԍ�/�fr^60��YN�~�J�\w��B���R���%�E�z"B�XlxVHYEB    fa00    2a40�>ԑ����9p0��z�b>/��$6�5 Y���"d��L�R��n��}�%bؼL���te�u�j�|���Ǹ9CJϣ|� Fz�\�d@� y�^
���\!��eYar��@���2�(���?�4�U�1?��o�����c�|E�R��3_�yP��R�_����O�_�bq�x�y��H!�R�i_�ݾȞ W3�Ɏ�g��yT��J�u�~*��q��;Y���o\Q��U
��Q���I���je�Z�/��1��cY����d��rn��
pb+v)M
�W{��sCq<?d�e�'�<n�ߩr��<�v���:B�,�XHO%L�NS?�]VP���B�Yf�}�0��R*זȏ�k.h��#h���it��폍.��p��^���yܚ}��Z	.��K�D��ܳJ	��@ݐ�}�`�<s����J��B zh��Y��Q�����]��֜� K+۸�Nq$�����3�]J*�a{ˮ=D� V����,���U�4S�)���S��H��9�D5�� պ��@����GA�#�6��ms��r�6U	v��~���'�+93c�"��>�r��� ��n��j�Pv.��f��QaOf靥t��
n�V���'�G����P�d����ׇJ��t���tz)��FjHQ�
+��w(�QH����K���oD$d��a�
��&��`G��l �$��,52r0�U-���8o'CY>�R��R�*"ض8�o��h��g2X��[��̬a]�v'8�'Y�l�z�|)�ɑ%��~|X{S*js�m.�3S�:t�	\l���Q[X��ȜIw�E\�S��e˷5M�!v��?�_L��8F�ӄ�f�F������(HX�$\����W�
jqQ%=�K0C�df�|�V��R.8q�C���{�����7CK�-x�s��U��|<����3nY�k��	��Y�,.�i�1.��x������*�5�����2�9v����*��J��d���o����'��Rb�=@N�O/[k/�� Ž�Ep��� 3(�l�����6�Z4�Z��[�K���B��e��ZK���<�,g��Z���H�A�
�i�2uۜL����=�1�����B�1"˹9���#�N���8��q�?�. ��t|��	L1c@U 
M�	:K�d D��'�]]��6��O/���LGcѫ��9Fֻo��CA�K ����ߡ�=z��4��0k��~��c�ɳW�J�2�>n�ۀ�^m*i̊+��u���D���u�iv#Cw�Az]y�.��O9��x���|%�G��*uǱ�N8��;v��_���F>�ߤ���U���KT��	j\E�����+�~^��.�s~L/�
_nɱPӐ'��ҵ�bev����d�Zin!��T/� ��˟	!'�׶ŴP��wץ��"���e���!�j,���V^E٪`�+=uS��yχ
�4��ݾ�=gfv&������ 饼��њ���J�Ͱ��w>8��zw�),��lch��$x��*n��+�H���7�<�_����%�.�ń�0�kA���uk�XŰc̺�m�*8a�[��Rq���H�Hʷ��L�^�}�T�p��'��6Ǯ�?��R�	glbp*�p�n��� B@op�T0Z�@e	}��Pߖ��=��2�LK�	���aE�٫�]�[��� u���<S�r~=���vb�	4���J�R(1�|���P�X��U���q����Z8J��ٿ���p)LK�KȪIߤ�c�����ea��ס@��0��~�_+�Jg�� 1�D�7$� �Č7l���3�M{Ȟ�/;̕����$�6���=~6���1�1�j_��u�������U�GD�-ɏ�N�,��~�p���N��/x���/�#��cdܟr�#����n���f�|�Z�{���gF���;�@��}쬁n��֚˭pv[tN%BH+pfu?�,�/6��`���>�-�)x�cEHltg�+s���2�$��>-�5�8�
��"ޭ�_��t)�g���z�
XO���	u��I��m��b�1��u=3#��o�j"Κ�[�M�j��#��i�o��+�K�okq� �QY�f������a���}΄�ur��Aq�y�q� ���A�!#����˨�n��כ�2�4B"~	v�d1�,��~�k���Ro�t�7�7�r;��TS���d)�2J��j�#[L�w������8g���S<puNU�V��8�f ��A.#��A��E����3���6XʳA
��I=���>�g`�>����]��H�E���*�y��G��_H� E�`�H��u�s�5K���ٕN�=`��nO���GF���;/��$bo���-�&k���Ѳ ��|j"%��D���E�x�s�x�������p�E�B}8 Z��CCjs��s�{@?�y����� N�S�y�lf/E{XE�~�6J@��p1.&�	��QRJdA*,�|ͤ��L�� �f��-n�s��dY��� 6Ϸqb�.�w�1#ucT�EoCz��@�h�'S����On�lq���MH��l~��З��1�I�-��a�ҿ�����Xfq9�L���m���������料��h��:�7�&����+5_��8�5%�S}�AXL�t��/5{ʶ��zX�WL��U���P��hq��{z#�Q�`D��9�)l=����+�A�D�Z���s�bF�-����ķ������v�X	!�9��¼�xe�?X��~|�`EGā�J�JY*�9��{7�� ��J⺲�v>q��S��|����j�Y=�x�WODo Kاw�W�(�U�ܴ��>8�}t��8'<�hB}����ӂ6�[lRW���I�=�Mf�10~.qȕ��
+,����h~�(�Zv���e}w�<5�RTŏ�*Ժ��I��0��!�D/�zM��+b�<�:Ì��|�F��v��qƤ�R3�Cy����L����n
�xT��EC?��Rp�N��ƛ�P}�V�f(DJ�~K�S����-Rw��,-�9m�ISIyc����ɘ>ܑ�/�8�N�
�v�(�i-��w��j��dH�F�.��f��f�!���h�\�C�;D���3[�'���D�V�ta,���Ȝ�r����5�uE��4�!n��.r�@�6F���ԱI{~ɼ>��q�%!u0�B�{�
c�s��u���[�����M|�ȯ��x�2�,=��7s��f����3SU�F"~���|pv��%��|��JH�_]e����QT�i[sK��Mveay�������m�(��?�� ��/�=�+1C�7H���a�"����B��Z��sa��'��C]4����nLu���Sb&s���
� �7�	�pǙZ�>2��A�;���R�_�1L\�b��������㓲�&޵�K��;
����9���hi~��"@������j���j�SM�T��0߳@aٛ9�y�^��F��1q#��mTpe�]����+'o��T��;�DU���oˇK�G��^���{�@����=$���B�CТ�����D�dJLd+�}	�\he"����z7ZY�<���;L�	Cn�"ӹ�)�3P������oi��H|E�C����1�X��\�IR�FC@:n�k�&{����W��ϖ��hi/g_vG��i]G`$�nT�)����n-G��YPC�/�IP�i�"� )0�ѿ�����%jbxnq�ߒ&���z�C*o��X���r��*�Q �T��6aT73A_��eov�td6(3(�%��%@g�� �Ҝ	ڢ�������.A�>F5ƀ|7�J���JMX��xy�x����
���񹬟�vxm3���|#�=��r�)�.��R�Nk�"^��qq����"�Ff���F��F������J��_|��� ؘr�]�{s�l8]�[:<ۘQ~�l��@�>�L��L}p�G�!�7^�86�z�M�k���Qo�{�u����A��pO:qF%B�P,��Us�M%�'Z?x�	����,���;J&�ա�����$"�CI�܂ ��OĒ6R����jȰ�����o�90��)�,q	��-@�0��F_u�ԟG)I��6����'|�!�8>F���,wdp�u��K�I�ou�9F�;]�Dt��,|=��p�&������n�l��30���.ݲ�`|�6�5�#*�I�����D4��R6������h���r���b-����*8:�Hz��)�D��lP���lC�P�]�K`3H��À
�l����XOy��T�x#p�dT ��}�{��x;����ʰ4���q�$;���\��	G��
R��L�ٶ�r(z�1�Ê>[�w�v�h�iL��cN	OйWT�D�#3C���S�R�.��\����Xh0f����BPR�Di�=�eKV�(u��5�6b���T�<ꥒCiRJ�eh�O���q_O�ΐMb[N�w�����_!t�jY=VJSd�Hѽm�X歯�rA��8�YABȪ���Ń^�J��]e���)���v����<h� ����$�#���?c���h)�&^?"RY6��/�{�˕�v>s�r�>�H���r=��i��G�GzZ�%���o��
����׃^z������\��(h)]e�(/�X�h�.� b���3 )��WZ'N����W�,J��-�=U���F(vL8����<�n8M�:Q~�?��;��6A�L5k�Z��n�<T,,�H��b�Npb���Sq�ji�`yv���:-qʱx�)j4�qNugz+��%խ�OkLck�2k�6�H��_�xg[�o�{��L�߱袘���w�/ٻ��.uB};���b.Xv��=�l�!��xۑ�ϵ,�t6ߚ��E�(�4�H�AQ��?�e�k�W;VM&�G�ɋ�ف��&)�`�J�|0�+� �
����FPJ���JhV2Q�O+�aw�N������#�G�P ���d߮�)M*�)dp����H����VA�~�O�X���c,��	p�J��S%��t@j�aO��|(�lCxŊz`��`�&�i��?#��B��ҁ!Z:�x� )�hK���N�Ip����e�AA���L��Ԕ�*<�F��m��iL�J��[[�,����K��$�5y'���"���҉����M-g ��#[O�~SW�"�&���S����N���H1�٨�up�d�O�C;���k��^�x�w���Y�E@��&o�ST52�'%k�fHTs?���*Hgl����Zt����f��K>r��=(���W�X_Mu�z�U(�=��u%�d1� ���]�����9�j��4���ϣR25�i�@h�̂o�p�$|]��M�<�VD\{'�c����)y���7�XIM�%�e�Px{�sdՋ癹2̀a(�q�9�w�P?��j����hgֶ/A��6L[/���7X��^O����e]�7���M�b����jK�P���YAE�-#]m���}�����V��"�΋��j	HV�����A6%UX����;����_-����31�8LkK� ��&PH�F��!��1�&c�У�O ]����w�J��y��ᅢ=;�Tt?�8�K�`{IO:AC����& g�0{D,�L笌)>����'L���Y��J6(�*o��
Bנ���v���o~���`O�]X@f�4Rz]X(v~��pj�9�k�rX���"���J�Pȩ�%�>��Օ���Ա�[Sh�+��%#*\!�HmJ��?`r�R�#��7'�<�f0��>pq���u����g�~*�E���C'415�j�?w{˽!�|qn*��Gf�!�.Q��T�E�D��J^6&"#P��_�3�3˵�N�@LmA�VT`���S����c�H�C����>ݱ]�W3�{E���0f��=g�6Ӵ�P �U���:�c-�3zî�0���?��`�G6o�%�����bGQ<V�T~�*VP�٩e΀�t�ˍ��_i����aɅ�&���7�L����[W��K'�^$�|x��������C����Rlw�?��x^O~��a����j�5FZ2I���>��l��`,�7,EvV<��ms��sw)Żv��۱�>��CX���XY��B�Y��ص=`������3���y�������>�ͤY�V'�3W���2�*��x���S*a.eh������_�~�#Ϝ�J?��e�+�`�<_Ƚ]�I�ă��g�������I7@�݃��V>��5�\m�{�&R���D���'=Ѿq�HXzb��5�؊w��F�Ȫ~\����]��&�Ϻ���+��=����ɪ��J��i��b�*�2��"�ݓ���qg(S���B[$�1��ِ�EC;T��Ua�éB����d>!��j�4�q��/�7k�c�����Ow0�3h��{6��p�RɄq-F$�k��,	�\��r\���l�T�_����o�hAm�7��Qe��LSe�����W;�B���:7��o��~��.�ojة��I<TsE�?
Ġ�Y&�u�S�^� ����\0�yMi3��:�p��I�'�O(���<�â�r�܇j����*H�R�ޘ�l�y>�5��rm8�B��W
�/���\hLd�iH�,FЭ�S��E �m�����hN	����8�z�Bk������|�J9\�Z���Sʍd��
��P��q�Pv�!̛��a��`����h�rё�z�}�R;c���ꌡj����+V�.�2��k�,��1�B�I�l|�R;������)j��HI,��u/5�z�8���e��2$&�2�F;��s[ԩm�7O��M? O�Y|,�WIG�&�p_r/��%�1�i�I����E`���!9p��4"�����pK� �"�aq'��_ !0��:�L	��O8e�kZ,QQL����'���TSC`F���7�J�^`���踤W<`�݁&^8�uۜ@�8n
KO��yz0YM��D�M%�ʝ��e��r���$�I��|�yn��uWʗd��ɠ�/'e"S	p�L�#j�^�
����$��P�bB#��4,���t8k�JgiS�ٽϐ=H'GL%w�N�K��r �k�t�jG.��|�f@au���&�hd'��yc�|��=*&$"_����,`I�e���{�IL=���ki�����;�$�K�Ȫ:��3�*�6'E:�#�C�-�˔7��9�v	9��;(	u{�r$�������[��I�xiiG��O�ܡr+�)b#���P� �h>y;V��AƗft�.�����[�нꍿƛ�IQ��$�*�����b��NZ�*�ж�M�j
/v�����JL25�=�M��p-�h��^�r��g�p *�X�i�X����>��P�t�L�GE��G��,9����>X���A�?Ns��na]D0m�6!���Xa)�t�1�,i�5�b4������1ٯ!Q�o3P"� ��z���V#├�����P[���"d�j+:'8�tzT��<<��%I����tT���ߓ`�A�G�\<:������=���p7G�Jj]�T9��d��d�s$k�*�*�B�K5�S��V�r�c��9�Oo���4�� A$���G�$�LL��\b͌ͽx)NʯG��͸��r�MQD��dX���Tn��^%h&$�a��>ߨ�	�Q7V�0�{,h��ز�謦���H����r5�P]g�P�ަ�Rgt���'l�za���L)J�l�<Oo/���ɺ�'b�P����=Q��a�j��w�f��:�����a '�����v�nS>��<,Q�]�͢��>P�K��~Te��a'��D87��<m
H������>��]���m�W]5�"G&�ۙK~�<�N|�������X��]�^?�[�2g� �p ���̌�~�th����� ���y��/�C�h�2�Y��_�'Gu��cp�"`�WSf�`�S++���ksR�m	���C�U_ѣe[*RK�6��H�Q�'4���	��vOl���L&˻���{��F:+9��s:�mQ�3Ȗ��l�-}�J���d
�9�z��d���.1��BL�#�F�B��:�җ����Mý��1����:�+i�(Z�d�b��=�j����j��W��^�õ�a¿��!b�Z?���;�P���uIˤ�L������t��&R%RW�؆Vr��!�v�`����Ӯ��o7ڝK9ql'=��l�����g͉n],��aN!��b���6�>�>�} ����*���*+)����v�/)���T���Ր+4sPo�Ż�:��z���v�����z��Pj�t����P���̷��p����U'�5��]������ ��t�r���{
�(򷛥�3�R�
��2R��Ul{\,�9+���]����� �d׎8�[�hE����{ŧlq������q�w� �4���ϫJ�Iyk� �e�|�W3T�!1`y�������~���௚��M�lRX�  ��Bye�Z$��l6�v\W&0�mt�J|�|/�-@��B^Q����@g� �(���j��B��]J��!�I��ó� &�	2��̿��n��ݶ5�P�C�J���ݥ壬W��p�Y��������gX;BՓj�bĥKR�5^})��������l� B��|�՟f<�ʪ��_�
�	�0��N�L�>��}��4�œ/�@a�4�q�/<��C@��;[=3)���mW����I���8�A���1�v�'/D�Q+̝P���Qn};��V�1>mN-���R3�@�c�48D�A����f�-
��yy��~w� �*�s1����go����ZeݮH�!���r}��{��v(�\۩��&�Mh9��:oT2��^?����Y%v���)fA��ڠ�"u������^�0�y�	���%���`�P3U<���0~�)��/�l�OQ�����1#ՌA����
!���Ș�ab�)�W1�֐.Wt���O΀V��a�4�f��m>9�/�հ>�K���S�7���}!�q����G�Ƌ��C�oD�#�ۅo���:ś�Ou�nG��U=Ӕ��uE�T�����D��Qa�Irݘb�9/�sك�P��t<�9h=�7�%�Fd�B��I��ω�/��f筧L�S�f;��ƌ�z
$u?Lzn���o�?N��nT^׊��D1������Y� gf�h�D n�Ӵ�'��Ŭ�����-��"�y{���.&nz]�-��u�ϩa���KPu��ݶ]��n��I��1�R)Y���	�6�{�$�=R,�
:V�@p�P��ݞ�h�H���<��j��Y����g ��=?̗ʥ�b���0�&d�@(�?r�vo�$��ağ(�l����f����Z���T�q!m90 ��!rr��<�DV�ؚt#�'��d�5���X�f)	]������/V"guS�1�ޱH�����[a��|��/Ju,������'4,m:c��ݳP�#Ű�lUX������Ŷo��vޖ���i�Gf����/�IyR���С������H����t�*���\��r��-A��fU�}R�
Y�08���*N2��y�{�q�=���I�3�|O�C�ߋM�#B���k��=n�<������H��^�t��Į�0;<*�W��Z�Lԥ��=賢��Du]�&鶎Yk��4M��c�d����83����r)�U�cfyύ�����p��o��ε�9���Bu��m�}Y�-�#�������P�0�VQ�j�z˛|��	hS��T�J^�on<'����H�)��r*��*]q c�&g&�.NUO�f'&�*޽�ކi�v3��s���L,�m����0�/C�C1 �;ϭ`�ɭ�ⲁGQ˷������i��#�5�N���O�3]���\g�y�U�R �̰��G��t�AWVLj��EG�Nf��nMߌ���G�3�y�}�(�7UG�VZN���r�$�?�=�h�K�`"7����e~7i�E�mI�B���E0�����⌽��w��&�,2̆�������ܔ'	�����[~���KS���Zz��3���1�"�[w��D
C��À��D�ar�Du+	~E�����¿, $�-��&�O*�4r���O=w��wz�A�'��.,^�7������w�(Q/�"#v�4�w95Ft��o~x�ZN�ՏI{
���	������GpE�t�=�;:#g4J����{T��U�����
�|�^�G��3P��ڵ}���L5nM�)'�n"v>jwUW\5=q|���TP�5�\���n��?vI*�R�*-W�Ѻ�S�6� �x�h����z���X���޻��1
VIK�t�qr_��)�F��M4�� ��+�.�H�7r����q�ȃ�|�N�Y�B���@�p�L궙"�!�R��]wh��6�^��Y62}��Ʃ��#�SpwVs���#��hP�lB�,����e�*�B�6�>�݊�G��%|�S�QT�ݚ�;��-��7�>}��
��?`��k�y�E���)|&� z�}
8�z�wr����� ����5.2�э#��k�1p�X�����r�����|XlxVHYEB    fa00     8e0YE:�����F�Yŵ���
�gb-	��F{zx�x`VK.�}��:��B	�<
9�0L�76��-,��ҷ^���ƴ��شD�P?_��>��,��܅#V����|�ǜ�k^�QJ�Ռ^:��C(#�:����[�E ��Y��K��&�R*0Q5�f���V�g9d����V�3��	��+��_cC�s��������W>�սN���c�<(�R5z�[�Q��,���հ.6�W�����?�gp�E��e���/���[�^'�"A|	�"_:b��k����:]�tP��9ĥ�:����lx�̘ͽ�̙�YҦ;b�Un�6�K��Wt :T;�Қ�]��Mk���Ki��}:^^��i�k��@&����QX�/��Ф5TV�	��l�D�}��_�C�1�Bvo����9G�
72����*��O{j,�Bb��$��j�J�n\��T�6�\:���C�<�as7�~��g�	��f��ȏ_�7F����%E��x�rը!|zs��FI?bn���%�s�%"��ݱ��Y�n�L~���k��4�1��;�'���\���V<r���;a�A')�'������A���~���6̉T�w8��#� �zj�ض��5�M��!(���5�_1a��.B�W:e1����O���(���Yʾ��Χ����-��4�v��$��ƪ��ʔT��r��{(��S�b�����C�Yv�~�	�@j��F�޿��w��t��}�$j �f�0n&{�!���rH�댍ȥJ�4�ܼ��ݬ,1'�_��H
�ϢƪW���D���)��z�:A�N3���v�PCw��Xf���O=�Y	*�~�Y;��V�ߌ���1�d�{6��!����F���셾W���'���3$y�<�+�5�zV��4�@ ��rc�Bl�
��$���YX�>k�����L�N��x?���,Qۮf��?c/�����@�CUVuΫ
�+���ː)ޜ���F�;�J6q�ǡ���ճL�z��Q�F�ۊq����y�]K.X����4f�n@�t��kdR[q�d_�MJ桓���)��R�$�����7`�B2��A�:�^C3�x��� �z)�����0�C,x����K,+�~�M1�RgE�FU�!E
��+�p�P�طC�˕�m�Q�:�Y 2q�TT����X����RC�����8X���`�y�������je�E�r2Z�RF��0Q�����Χ��2�h>b.r�F��ޓ`�@�F_��K��j�'�=ޚ�pf;�A�!��ɋ+�(�K��*�Z؁C�0DD�>�$3B�:�vn�y(��Bz���ma	$'�r�{B�����������?��|�"����R����׏ή�	ucʾ�v(��.>�=�K�������G!\��9����*��S������4H0ί'C�b�ͥn����0XoFI�������:6����o �p0D��T�Ӣ�N�hj��>!3���~=��/κY��c�U���c
����xe� ��i��M�����p_��=_�3�|}8 �l� ��NFRNy��B�H�A�AĠ2ֆ��+��e����~��h�H�PΦ�|+p\��½���t������54[LQ���#_�I�@8�'G����	 ϭ.�W����_�C�%g�����Qm
Q D�}�*|/����|�x��F�\���z�7V�6���)x���=\��E�ј"BZ[�De'!/�Օ\)-�]��N?��E�MU�`9*�%�V�&��s6�T��L��!͆��8Hà��I�ĝ�9 ��<݀K��^�{��*�3�6���b�H�aslv��T�u1B��_���NӋ�.{���M(]vЬO�l�c�E���i�MOMl7۾�֦ҤbP�c�	P�1�@�l�\����҂t��2�MP��c*)����.�O���h�����ԋ��~3�pFG�5�k�ʽ?�oV��(+���i�.�)��!��u�]��������
kyY�d������29��qsQ���h�v��։B��r�M���:�Q�h�J٩p�c��J�U����W��Q��H�:�C��Ϭ��2-�uwP�b��.Sh�2 ��c���C۵ߢ���s���؆�뙞�R�5���N�u��^^�E$X�Ai��F8�ď�TF뻖`JR6�`��b���#��J�&�ۯAw���w�Gڇ�әBq{w4S}β�dO��6�ݜ܅�����rsXlxVHYEB    fa00    1110U<"�"W�	��O�e�lR���h3ђ�H)�ɩڐ	�V.Lsx� ��>��v�?I{�ё�]?R	{g#�J�g�ܦy(���Q�J��e����I�J1�>�k�w�ye
Y ~�g�=?���^��/�MU�1���B��|{���A{�S�ug��rᓠSr���5�^t�q(`�T�&��]<=at��gH�+Cw9l����+�[���r�Z"�m������`z��E���lH�3�]2����m�������wO��d@:���aR+�=+�	G��_p5'��!�����L�8����c����k���&�9ȪZf��*�������D��(�NC&Cf��JR�-��o�x֩p$웩Z�؄w�����JO4�T�q�d_\��nJ�(��ˀ˙�#uV{�Nح��Y����#�>~�ބ%�v���JjՠO�8�\]���+#��$%ȼ5�~��A�Ϝ�����W�Sb�e���8�>���ڛ���7�զ��R�����j����8qibƠ�i�2e8A�%D�^I]��G�k󪳄��������tT@���@������缟(���yRA�5�����Ƈ3�s�3�T�:��*�3v��t���jg��I��L@��~��H|�i:�Gn��7��ܿqCv��θ��q��ǜ(귤C��=A�`CD��TAnE�6�v�,e� g
TJ��ւa^�\ �߆JY��R���������u�\�	���̽%��9?�x��(g���J��f_ꊔ<���a��	�F>9 r�С�3FrH߿��ˠ��AK���n���)��ǅeza��\]u� HS?�^���Zp�vg�;ލ7�y���C+�}z�r�>�Wd��W;=^��nUR\b>�0�Uq@U��񂙘���%�u�uE��;с�[Ȃ����5V�A¤��f�a!湘[[�Ӡ	�|l�G�C]��a^��}�5�MY��w �H�A�+<�άz(��PM�����k�'^FN���I�|�P9�	���>�D�T*5���D!�௢*٦`0s��N�`��~Dml�~��}iAX��	�3���;��VbR$p;��\^�gCX�Bn��y+��B�]v�� ������V�0m$�.t���L�K����~�/�gRHy��מ��󾛐����5A݌�!8#:Jyn��X�\��.�$Y��۷�Hk#��%l��=�<��C�#��j@~��1ky�����E���y��f1�._i%����o��{���J�������ֹ�N�\̃���H��H����+{'[�e~�矞*kB�XxB����&"�8�\~��~t-���Z��m�����5UBX���3�}2�F,�x���#IJ��`_m��8!�w������D��W���C��e��`+��&�(���Z���vdHR!|���)Q�C��H_zi��cHOY���d��N�����$�D��c�E��b��m��b'b~�c�)���\to\��G���!/з��|4��v�2wt.C|4qL��q}6�MyM�4�	�?��-�Ul
&50�&�yi�G���Z���/��Z�X���R\��(V��}N�ls�Ӫ�Pc���2y�\��D���7�0o:�{�Rd�u���U�Vi�L���.�}����0�K=`)E
�����>B~��)x�S����1���y��#U�Ȯ��99�'�O%���v�.�߽vY�*2��A<�����U��,)h/��G\u�!y@!�!ȶ��Z;T|h?���8ˣq�F( �ŗ������r�y�.?���x�J���3��9���,��G���02���
m���-����z3�o�E?�ˤ �S�@:R$��P�����1�NLFA!5J)q�;���ȚY���)Е:A��rď@9uj%��殮�<)��4�+U��֯5q�HT�r�d�� [o�����Sųg_~\��o� nRqCP�FLx� ��@�t��_6��
�eYA�v�\�-�hg0n�k���Ki&\�%I���Y �9����9�g&G�b݃AV��U�4����M�.���}�J��af�DD��6(�>G`J���|�����c�a���H`C��g7�̅�!�������1R0%��.�ty�b)x���d��">����Ֆp�z^E��>����@��w��P#��8�o�pm?����g=�H&��"��6��-�g�YN��l'�Y�����#�?o��>L�aͮ�_��ܟulяWǾ�S߉�p�K���d�HHS���|��u<�(C�q��>~�p$�P��_�C�%�@}O��%ú��Pzw�_�&B�w&v���S��o���z_S�����sDdG�^(� E�sKݎCVճ��^�;��d�PV���Ϫ�B#�r^��8��:ȄR/0,��վo*YX��F�U���|X��</�r���
J��ʲ��@�q$�M�N�|�N�Z!X'��<��&�;
yx�gV�E7�^�y��(ASƜZ�����,��zr�w�|<Ÿ���-����U8�$���uL�@ָ)jӽ��1/t������ݎTcˠ�cc��Y���>�s�s^�����kN �c���i?��I�h����c�U���>�с�S4#@�O7e���"e.e�܊�$�v�C��4�ko_�wq_�u�0��>�P����)ۣ���)_��ߥad�Q���i��{29�Dk]<u�"<��3�A�{���@�1D��ɋ�~�pw�x��\O��,N�m
�[�#�f�D`��j�]�/[E� �,��`pN�zg]�����~L�>��zB����u�wx_��57A%$�_�M���@6�����f̑�`��u����N!��9Mh�R�%��ҽ�k*L�B�PoE���fҒ�O9�܊�V��tFQ���f�ԍ2w�6ne4UV��HJM�9F�{h�ɶ\Kau��580sg�D�+�-�l��{-���H���T�9���rے<�=A�8��xSƎ��6�!����&��ۻ��ȶ6+a�;88����R�����SCB�+���x�"2>�"WE�N.C�j����>�bپ�<�<#ߪ�w|@���6��J�L��<����IR���r�K��n!�lh�<7K�&Z��3��.�I�H��MSD��@�������~�&�uE�z�.|ڢq��;�:�ݣ��I�
�z�X�T�T�	�K9cF:|%�F����OSPQ%�0����`N_�t�]_�N[��~<��7�������x����\�k���d���:[�1U�5��u�^n����5����	F�䵏��J>R���ug�
�g�]ԾL�*��r��t�A]D�M����;�Y���L��Y��}��.�~�FQ�M����+�j�]�qC������C;��1����8Ju��h�l9�y�w�88��\�`�x
/�����I|ӗ*iY���C�\'�~ �j\o�L�-�:�[%r}�\�P;Q?Zkm�]U��mT���6oiU�+�����)�7y{=���o9x���ed���+���s�r���e�t��;��fK WM�^��5�T8:�����*���,�L;���`�0��xe�YO+�,���D�W��L���%zI�ES)>y������{hq:)[^�܃��u�U��(4L�.����}9�]R�𝏆XG��h$��ϒks�o7�}�+㭎�ut4t����Q+��U�63��Č�	�#r+�@��M�F)��j�9#�KYVK���7�O%���ʅ����r�|WȘrH��X2@��q�O� ��ޮZ5r�^��y��s
�Kvlܜ�hbќG(k�
a�oݫf<�9*��P��G�^�.Ź<�8�gtcϟVhtg��|�Mv�`�3�Y��;��H�?`Ci�u�Sp�h�"�_�,J��!�<�gJM�A.����O��x� `sg����6�~4�4�pG3��Y;Jh���ߖ���S��q�R3!���ٗUrIm=��9��"�(Uԛ��L	�I�H)��b.�wAg��Oz�DPU�d��T`m�T�G+�(`�4,�1E[i�\�{P�M�jJ�
#�͢Y�!��ĸb]چ��܍X�Vx�p^̲���r��r3�#D�_AeӦ\e,�r������ƆeM̗H�p� Y��Ex���P�bb��B��;��Nj�ZC��x��>�I3`8���T?Um��_5��g
��~JF�RM�#%���oP��Y+8K���%���p]��Bق��0���=�dOZ���XlxVHYEB    fa00     ca0�3*��{f��8a��z��g��`W�d+��j{��ɵl��)���t��D[" WZ�LS�`~��]�%�'}��[I���uWPN,"�q�ѐWv$���ySBv0�q��>��X�NmW��I6r<os��
�4�q�ӣ����y��:��C����&�e.d�.�����ĝ��.+&�8A��M��woz>_��|�m���ug�QF��PXkwH�e�a����4eUG���\��4�>i��G��S q#��s���y�N�B�g�֩�~P�oˢ��k�n�5Ƨ��� �Uk��6o���q�O�,����+8S@��8�hC�'��
���p��䪃�"��st+OZ�(Hiw�10��c�te�r&�o[��d��0;JD&���e �0:�3ػ�)���.*}�0VC4�Acu�����cʄ9Lp%9u��D=`�Uܖ@�Z�����?�x�G��i�Y��˳�6��Jg��]y�xD��E��c%M�U���0�Jɞ��L�f��X�u���藵�ϩ����Z�o�,Ɏ�T��1}#Mnj�n��Ze�p�X�xϕ}��u���a��Z�Y��xt�U�)q���ݼ�K�����\�k�����-��븩�Ovs���䠬w�Rҕe���CW��zݧ˂�I�Ҍ�Oh²�CB0����X��?�W̲���u|�o�򏯾�zD����+`�'y���1h�_ܦltU6j��_Sd�y���Et�T�rYr-He>�<M��� {謳�k�iR�����E��<ޛg��d=t���5�t�}�u+�XIƹ泍�ѭ��V�
�i�	F��P�H}����I_���씊�m&@:�A�E�e��{ԛ@p��C�޷^��J]*3ߵ��^��V� ��#:�\̢�n¥淨xP� k�����[7O���T�0�2<e����lW>z�xDC��>,<D��������W��hm�a����y�����BZ|���? 1�1{���ӌ��o�o|�z{���P�>�Pf���'c���|Q�JG�6/��v{oH*���c:�]j�/���N;���F��o��3������]���]b@��q�K��_&E��]3 �^����_{����j%휣��
HP5܉vLm��~���؟L�|��j���T,?T.˨T���6�����s@(����#½�o�|�I'�����h4�uV߻R�/g��E&����ae��Zf�r���O������Sӏ�l�����)�M�%Ҟk��ˇ	�. @Z������UZhO�~.�U�I�>'㹤���J<iFƕ�TjM�p,���T�e��"R����@|2-d���瀚-e��A&"i4V���C=��e]�)����*��
ԇ�et��n4�;����7��>k2y+D�N6�N��SDG[�0[��A�`�D�wǻ��vS;�b��\��k�C�S2/�EvɁ��a�^ݩ�c����H�e{��*�I�}v���d-��%�4G�}a�]]���:�N[PK���O�҄@%�^�m��n�p<�牉�CrWIc�^ք���}��
Z	�N��y��dw)c����s�aɑ)m�\c���M��}��+$��Z�.�	�G�>r���y��~+y��Fݡ��>�f�n��2�ʐ�qX�y09Dڶ_�⮾��K~)�kʙ��n�U���(��n��k�����b/�q)�b���WK�,����r5e���4����������Ҁ�� ��D&-[����i[����B�|k�$�{a��ĥ�2zi��������h�z�$�u��1Y���[����޹w����Xx�i�IQq��0~�~zxZ�J$n���U����d�X�����C��73��tO%2��	J��7.�ov^�V2�R)�A�'���R�<��s�8��X;B���C�젉�]�u��j8��`��I�h�i�%�1(���G_���i�j��m{�xZ�qP�� @َ�_���RI��5ق�7mA�+( ������x�S˫����jV�c/'q]����T�K�'��'�Ëp/E�}�r� �&����9��2v���9	7o��a�?�>�E�T��%|+�~%k�Ч����1J�'�_�(�g�u��hʽ��?���Ϙ~bUŉ�k�7�]�'����V|�ے�
���G(m�6����x�}Ǽ]�B�ܴJSQañ�%�_FI
�c�#\��(~���B�w8�L\����Wc����S�L��g�t��|Dpx��1�)9e��S�)n��J˃�d�9��B����i���#Nr!4��)1��|Rş׭��(g�qb��U��3.`D��$�̾�YjA
�A���#aA��6�5�W��p!�����wc�{�瀉֎��{D�9�J���(���V����}TjZ��PU+%�v(J���,�ׄ�&�}׉(�!��NRlqG8���z�ǂ�I�Qmf��7s��;���x�P���"*Q�2�`�ar��2���e�i���`މ�r����q1��'�#I��jVZ��ԡ𾽾��@fJI��
���]����20�:�|��ֻ-�Qt��e����+�<�ŇS��a0]�� �>W�a����,��N1�j	U�0[5���b��.w�l�R�J{�u�TM=W�j��1�?���sE��D�#<v�F�?����<Ή'���-�u��mB�o%����Ο����]�Z����D��4c�oj�w�xt%���qa�̽|�ߊ���7DI'D����TTwz���l�v��Ru�^-�?��˧Y=�`�z�4�A��C,)�y�
el�%`��F.kvL$SX����֜�������1토���x�;$*Mug�\�u���e}lVr0����Z[�3;��+���YHهRE ���dW��#�B�D���� �'Pq�vn��[#Kؖ@�\]��@�l^~�.�J��|��?��A�
`�r��5Ӊ���$��1�@�g^M��<sX-A:�����׍NE�QY9��k"�i�=~d�S.��$��-zF ��0F�G��.��X��#4j�8�r������b=9�9�:����-W#&�݋�^�%�Vd���n����v��ㄤqpl�����%.Ew|k�"@���~^(�^w�o�#���g)켬vܟ��~/ʭ�XlxVHYEB    fa00     3f0�n�6��(�6��W�O�����h�,s/Dar* Ϧ�ߓv��W0��>�� �@�7�$,��wqI�� ���]��1��`�VL�9��7�p,���+�'h1���3+�5�2�)h�!?ϭǚ[�s׀5�)�W�'(z�G���.�����:�Sυ۩�t&b�+���r�R(�X?T�"F��ݫ�K����Ѷ�V5*���V��&�6�Z,Olp��Tj��R�`}��nL&�)���9�L41�ڻu	�!9UX���qf�R�����ٕ���P�wI�(3pLX��?�T�PRf4�-��:YP�EƵ�aG�)��#��n��6���!zQp�2�5`����xE��-~X�#���b(�x�W�S���C%P�D���6�����k2��+}1����$�֍䓇\'�'�^T+��;+��ӕ �`	dw������V���O�H1��F�"G`v3�i��K�,Z6wp{ej�!���@��:���92���s�|���U�z/峒O���R��Kw�a��4�G6�ل���7�R�!T����:���'�"A�}��ι2U-���[ݥIC�g�OA�㫀�G֗�F������Wp�x�_��&	^S�h��$���d���XY��g�[��7�Eq�ɿ��˳nIp܆Ng���l%:����a޷���8nP'/acENu������'��RC_ޚ�H�Ϭ� 3�Pr����E�86O.(���Bo�t��o;0,�7ѯT�3�E3�HK�ڠAt������x�������� wK�on�X�ǽ��k5ǻw��Q��P���x����hr�{R����df�\�ZͿ�8�tZ��.@th�c��Sn�t�̻�����b�Ɓ'R�K<�Ƙ��t#8���o(�~���#����� �����HAu��Qs����^��0R^��I}<L���<)V<����%L�n�����\Q0�v�yyg�s��q�Q_�ϋ�6��j�H�Z���y߂XlxVHYEB    8096     b20����w�L���v>n]�l6��y�[�8@K�r))%`��t��}�,�.�W�?pAd$�7Jv_��ov[�;�����uN���ϻ������؃�%����R�|�0,�NId$�E@rr|T���`lQ�>�"���V@j��L|�O­�3V��C���Fg�H������Ȯf�:�z�~�D��������
S��& �_�Ǎ��@��(/�Tn%7�&�6e�	�粞��<�!7X�;V�=��!�z����&���\��i�ĝ|��䮥N�ku�����bs�E�V=��`_�[��/��F�������4�zך��᢮�?���*cY�.c���`#�XS�܈F����$�yΜ ڞ���O�p�{L]-��EE@j~˲m�ǵ�tj:&��̚ �!_ (�3e �����/I;��[��b�MX%�-���Xҕ,�h<�ٔ񘄗�<��	Y�3��Ά�.�\�mea�ZMh�P�%����N��K't���fT��u�I�g�'{�]\��!�n����:A�%�M��7+���c�&���kVE�{��,Y���5����W�+�ɉ���Y�q\�����9����0�q��I��x�c�Uf��y�QS�W��q\p�ړL��k�2m2L_��zm�F�b�-������1��f������ �L�*&+���B�����<_prq���<��?-�ƃW`6i��F����5��R臻��r_��Q�أ���� ��?D:g�y�3'J����{���.� 
#�MFq|^'ݦ�Mݼ����;��Q�H2��8�豇�+��^�0}hH��{��ś���k�2m���ԠXB�;#c�Ȅc�q�i+�plC#d��gQ��Ň�;ߜ�����ۣ>�������xס| {@���T��o��j�2�IsZb�Z�ɂ�>��#U�5ă���M�C�ZW�窏�=��Ś�)�^yx�S39a":Lw�4~I'eh�:q\��=L6�^�K�1Hg#YEn����&���#H�����ܲ�>�l�M��$�����P�v�W$�2r�N�)�����C����O!��_@�W��oy3�ks�����}�Iz�/��&��~��HH�c��V����Њ�����NC������ق��^W_�"\�ib��HK��¸�j]��=��4l��4v��(�7�gL����2
��Q8~!r})�0w���U�������  �]~��C��_5��Ʌ���>Y35�@�y��a��K������J~M��v���4(bY6����D/����S�BF� �M@�r�3:�H�庳��A��ٺ�b��Pu�<m� �YǦ���~����o^֨��^~G{T6&����o���wB�������R�Gqq�{���~xҢ�-~j˨��N�rS��;��B?7�]A�<6�7?�x.E���9�~��#�CS���Q�g{�'E���u�j��\h��=���OUR�4��K\q	>��vG��)]D5�� ^���.E+4܃*���u�!�Q� ��^�&�e������4�𩇋(��aC/�#�s���5�}�Qu��s
\С{n�3U�Zot�}�.���6���ςف&��U��X*3�YvM��`p/I�d@%���y���f<�okl�Odl�w�����fu7�S�PTF��D�gY�|���i�<
���j�V�X����}���sor�br�^�c�ĥe� H'\��c��B5�"J����#w��i���|(AW0B1�tچ�wʢP�����y�0���2w�ҠQ�?�u\:	ʽPYj�˭x�	L#h�r5��V�d��i��D`�c�\�c�Z �Y��I�����~��:�E�����\�x~S�%Y��un���l]<�/���m�!����B�=��	3��I��D�/\%?��,BT��-`kJ��דvmR�)���u<�u{GzI�{,��b���p�đ�"�@)`[��1����*n�!������:�M> �ߩ�����6y3Χ���>5��5��`�Q�V�n;��h���!�׍AGr�cf��#�7�:����d���0)�=6�̮Vd���WǦ�2��z_f�@����.&���ZT�9�LW�į���aEѣh�Ld�c�<��Z�����О�"*����b��L�[ -05)M*z�~�ŗ��]��ghKƄ�m!٫�B��Z��oʽ�3��ثO�@)�O<��������S�ި�P0��z��s��yR|��<b�Wkђ<!��bGd����4Ӆa4���-�6��w����Á���<aR���);����`2�%$EZ�@\b�����ӿ@d��=_L�
��rإ;k�Ѱ�A�(@��;�D6mb�]�WW�sեGLr՜=��혏"��ߒf�ٽ�s�z����ԑG��i�8\�,��0p�Ō�q�up#�x�	���8j\N�+TR��^uY	 ���'T���:(%{w�B��g����KFƄ���4���3�6�MDT��P�9�5��]�"n�F�zO��-}��Y)tU�� ����et5r�	(�<T�������5"Vן���L�Y�$Ɇ���0�BeJ�2I�lto�Y�R���I��9��8�C1�V߁���Dw������L+�����t�^�z׈q{�{�O�ɓ��8P�
V)w�%6e]����f�������CQ뜈r>r��^Q/"c?�X����C����"&��`�<> {�)���x�ǁ�n�1�+{쇓����s