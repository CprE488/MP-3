XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��*a�w���\C�"��g)��ۤ�BV�_�a D8|�]D�R�+a�]h�@�n�2G�+��I+��.73cLw_������\Nm\�~~w�8��.�uP�<�*�_�8G�F���6e�.�i�x�-�u_R�z��l�4�E#���{)C٥��5ݹdu���v ש]��
4�j6}�M2��)�������;���*p�b0qF����a�_'ؒ14
�>��3t�k烁4$�tnɁ`��}�2L�����c�Hg�Y"�ݗ�k����������g`�9�b��X|d�y�z����y�l���lh� ��ÚN�f�X��<� [���d��Tp���Gc���h}�-�L
�b~	�{_Ŝ��6ch���b�D��IW���f^%���J��}��M|H�M���sr>h>��}�#.�m����١�N���b�N�OU�����FM�w��Q|i��x�ǈᎏ5Ō����N�K�p���t EA����9��<4ߢ"�]쭯����xJe`�MO]�2w�F�aƨϸ�q�r��~ϴ��O`�p�&k�il�e��}���D�+}����텆&�F��j����"~xi�	����f����a�uu���+��Xm���Џ�"�ٚ?d�b���VdyF�r^Da P-�AC$�������n�zN�^�[6��?|��2l6����ŷ�)���T�=HY�¥m����ǫ"���?�l-��0�
X1�2õb�m�������-�ǭ�tzȴ��XlxVHYEB    290e     af0|
MO��Otl5��WW,�_�괽Us�W�R2O���fa�/���&�#��0�ʃ��O�hMK+D���R ��my�b;��s�_;���BN�#j��}�Ϭ�nl���g
i� @/8.��F`�w7;X�z{��l��&��zE_�~��I�βqg���g�P|R=���I�W��RrhGZ��_ä�:2�3_):����(U\�evOP�)���T�G�D�w�u2Pč{�q����0w���{�-7���q2e�VeKm�h�@�n��+X�H�Ŗ�,Ⱥ1I������gW>�eW2a}�|֢ ZC\�]����mW��m�����Fk�h �iGܑ�?�ǅ�>�O5g�!v9�<���?��:JX
�ԉRM.p��&���< ��Ċ~�ۘݍQq*h�yT|� �+��*�냧`D�ˑ���wI�N�ʐ�����-�����f!�	�� ��B�����j}[� �[b�$K
��jq(�$���ň�[����\��k�O��X���H9��	�L�q������|�L��}m��}���
"Csj��-��|�Ԍ�"�11X�7�Ĩ?��X��w���t�2�Sm�w�ФW�evܬ�5�#�R��	 ͳ[2n7���� UQ�A����~+�ƚ ��q��@�l��������4j,N�����
�_�x��?�����	�3�Z�.�'��CK�����dw�L��m��v�2#-��o��^����cZS����g�݃@A2cS�����op�e����MY���C�.
Mܠ�kJ�;rS�,~��ETz�I���������?���>�$�/�c!Ue3iW��S"~'m�od�C[6���=��֜�������e�Zz8��jُy��d\�M��<��-Yq/k��f��L�E:߈�W,;���l�j ��؊�I�(0��.��Ψ�
H�:eA����������Cq /Z����m �O^߿������a��@]Y�7�єm�P2�H�=�R\�Ẅ_yapE��Bz���7'�p�"�;dtb�)��%&H�-a��i��$.�i2+(�CJa6ޢv%f�Zg�}Z��u�`��`nK��9p�vE�	ɺA:`����J͜i!�%>*��0��T�@s��
��Nq�n(�,�3,Ҹa��d���e^��c#�۽�b�V~��NIv~��-7����q�iI���o% �������j�􂐚.Xu+\���oJ���̈́p��b��u6�������av��l<7�1�N��l�nԄu?=�c�h�	w�*I�X�j���{cI �O[|x�*�X�KGs
�=�oz.�y����d��/'r{������H��b鏂Y�*kG���g�#~�:Y)�2[_B������F�/�>
�k�M��lD�(���|I��d�\ctlԏS,�ke)���s���}��c��^V��ߣ��`���ݻBjİ����+2|H����9i�6�3e��=�������A�#o:L� �8���CZw�w�ZdtsY�|A�NDʏ���=ŏ�g�%!���������Ki�97T+
5҅��J.�8qr��y��~ �ÕY(f��զ��>���Jnߡ�ϴ�WG��s�0��
I���lp�p�U�j�����ާ!
U_9�
N��+BK&�Jn�<k�%[0�9c��(,�~ٙq=�sH�$7L��Y�g��gI��>ֿ��Yl;������U��Y>��-���L����*�?<,���>-��������� p)R'XsA�P�E���+���!Z�{Z R��M}�	�+�/�r�\F��
�a�j�����{�GD�U��pJ�hEd��>�y0�UN�)�-ضY�e��<�̴��VA'�ṭ�Rq���yc�Tx2��4�T���0����LȲ�^�ٜ���df1����٧�c����T��${�Ei�
���<��K��H�����Y�r9I\riSk�2^�c��V�IG'�
�`��77v͈�Ig�Jvz6�$ ������bu�>�P�Z�9���*F
@���ex����!���(Gw	x\��rA�᭰���gh:u�|;`���%�A�[h7���p�D�0qslȕw%��_��PW��j�@es�]�\�6C[ͱlr3c�cBs�)�KiY�P"�������:�c7
�V�=��^y�1x�9e���gm����H9�WN~H��v��=�$Fב8~]����gn��!��lA��4c@�d��8:��c�;z�~���n��xh��L���;�C؛I�<xi���"E ���y�S+Ӓ��h��
`x��R��J���V)� ^�����-�C]�A0C�̎[S�f)���������5^`I�*a���Th=�:�h�=: �U��?�$��а)�N��&��C��B���C:��)�������B�n<_9��P �%��h��	9h㕛���䶪�$?�5Q��7z�?�~X��%A
 N�D�l��Kk�°��ͫk�n�.�
���p�a�`�Ž����kߵ!"�r����K�lW�w��/��8���"'I&'-4��G�uj��U����E��:�92�Xާ��e뒄�#�`Q��� ��H�qI+4L�fM@6/1�$Nirx@�Go��+I��&�S*	NG��C�w�ƈs��X����@� �)]�
o%�?s���
=�y�9�@<���g��0�'��̽�m��������S�"�l��X䋸P֖�-2�����uI!4�����Hه���