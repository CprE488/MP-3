XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���[��h^�W�7%�����"�]�l~}�	�rL:KS���t깚��`�3K[T�pr��t��A���vq��2�������1��o�ʢQ^��UG8�ֶu��rz8X��e��VW� �����}� -\�-���>e�;�����
�_{�,��S��R�;\#Nd����^ǝ���Y�{��5��{�䓈�<a��1kn�`��^I�A2��B+���$��0�X�gB�Gq!*�������r#OV�p��2G3nDUe��"D%k��blL�#��A�	�9�Z!q
~���&��-#�A�S�.q�o]�0L9��(
�I��ŝ���t̄��k'V#��D�V7�i��Ι[c ��g$��@ǽO�Ào��L/�=�O�;�5�� �"�_�����D\��L3��䱫��=�{Pk'P2+3Æ��k�o9u��WK�Po��w*l�Xzz���h ���+D��],���;^��1���; WB�P�G��gş�{~縰��>\D�3R�3��dG��,�� �t"�lŝ���?�`��ɓ�!
(��a�S�y��g���$�In	���f@�O�?E=o�m��J���z�No��u3�.��h�ej+�`��)J�_{������#��°?q��vy.147��P@��0�b�p�))�?X�)N�b���"B��2�~[>M@k�#�[�{23 �}�����x�ԃ��F����e�'�SE(]Gp�d;*x�J�w
��Q9XlxVHYEB    4284    1110[�n?��ДN��P�=М�v�6�؃٧�8�������3�!z�?%/2mHgriu�F}�j�{��]. ���I�)y;��t�R��bG�9�Vݜ5�q�����f��>V���ŷ��
���V.�k>�;&H�O����3˱`o�હ�1�ޚt�Q�6�p��X[,IM�@��_A䐩_=P�I7<�=^��=�������P�+��;��c�)�L��� �-�ڤ�W��R̸��iÖ���1�b�#�(�k�MF=j�H��L�[��J�"լ|���,e+5��=B���О�0e���Fu��ngn�@��[oz��re�]mQs=zB���&��g9Ct�}`�^�'U�����f� �&�"�i��L�<J*�?�W�J�5�,�>5k�]��6F�.>�m)}oBEUO�`��n�)2�'N1�m�A嫜~4}�a��r��,�О�͈��>�3ӂ�DX1q��	!��2��/B39��oU�R;n�*�*���Mm%b�98�mΞ�Y�;�IƁ���K[��KGn^��������������\��&�$�c6��-�<����-�u�/n����Ԋ�1���������j��|?�R��9	`=�鋕��U�=&,��I`��L��f����(�ǌޮsr���&�����yq��+폂^@� ���}c��Ŗq��'�d.2F�������F J�Z�z����_"��6B$h��ea��d�,K�W��1�����&�/�]_'-)�r�(^�)�#,#����d�<ߘ+���V�$L+~f��M�&��g��y x�O��IM�+D��nC�qKg�O$����+f��zCӄ�������1c���S[���ퟝ����WH�|5kx݉�;��X��:� ���T��JZx�n!tj*D����~)�cX��r��t� z�oX��T�SiJd�P� /̼6=�E7�Y.�� 3Ԡ1��l��:��3r�o-���/:֐g�t<����c8�q{�`΃s�W��z�K���ɐo�I���W���a�{�Q*Y_:�}[���{iL�+e+<�Gs��d���MM^����89�C-���p��1m)7�-�g�|���l\�X�||gb�|Uq���<ro�+ux[b�}�h��
\=Hn���A1�u9��{��:�㟇CYl�.ک��1h�t��:��g����AH�0��f{ϸR�@��',��Gt�UK=~V��A�1��oU���/lZ���V��&a�g@�3à��-&$� (R��	?��v;h:<�$�A�f(�'��W��i%f1�P �}��䚭�b�\������"�zK���Q����d�D��uA�S�0#��~߯�B�+n�Q�̿ZP;�R��ƀ�MIcl�\�]ic8G�yiʼb�T`咶<���ᨨ�P�5G��|���gWșTc>�{���s䢽�;�؉�GE_7����u�=@j�+>��
��u���w$^�Ϯ)����,����	^6o`���U-dD���.�|*��D�<�V�gh��3�znI��+Z|��!��ߌ�0	~='�`�#b���7��~ј�5�^�51H�T���{R�X�*�)s3JEH� �D/��P���t�A뽵@Cg[�r�ǫ��H߷���:�u;^hz�d��pu�p�n��(I�Q��4�z�m��j7�\ź���*��R�l����x=��g���̺cc:g��VDV��ؘ�,�^G�8��(��Z��&�S>M!���z�C�2X�I�K*l,�	p^iX�4n���#��FNW/6�`)	���*�;�2���6?γ�f� �p!,����f�����(kfI��{����dthI�ï
{�Y%� ���r��e?���qĲ)\K�S�=O�1��sd	��j��j_S���&�������$���~��9���;�� ���U�+�,��dOk�%	��?m�R�����k�������׏���>���Vl��H�4C���|���*#�6eM�{oh���;�G�=��847�=Nj��i�%i�R��|m���\��Ŵ�uEr���ūs�R����١���;��_�RL�c�_<��M�h�\()��Oz��Tgh�ZTȻHq>!
�,!}8�U�B�^�+�	i�Sq�2�D{�d,��,���`��K`Q��� [Y1a���4l� �O��nDf����h�
:�+�����i�u����kk�4��xкӎ�G��%fy�PtĲI�6�M�#?P	��۾r~�u�"�ϯv�x�t���,Q�.�<����)�8ol?�7G��`���ȶ�KU~[�6Z<mU��j��"���A��^�,����L�-��̾��ӱU�fkpE%W�ݢ���l*TN��pe������bB�IR�w<��d��7�5{��w�ߎ.����)dz�ݟc[����6�o1n�U,���D�/�ʋ�ǠI��tM	A��F6��n,r/\�5�j� ����tsl�/OXj����XT�YX[[�#6Uz8P:�o��f�ł^|08h4\��U<�jm��m�(�$�Ie[�Shcx@V@ǋq��M��ma���<���&�Җ����c���>���aH�(y�m�[���4c��STr����C����#�J��������f����/�'���ᗃj+ۼܬ���}�6÷�،���ڪs��x~�uz�� >������5�/Y�mk�+W`))�����?�V�W����M_ǣ��z�a;y�߽	�a7���kμ�VK�!%;v��k�`=�fd��u����I����^�����Z�v߬٦��I�����~�>,�*qʂ��By��+F�4!����(�$��a��ʯt���>�$�3V�<Q:d+%6˳��ub��*��lA=~�,G	g$ ;+�3�e��z��P�r����a��I��m��,��_��#?����(v�՜$cf(����8���O�S��4�-���ð6��\
Nct�F9j��q�1�_K/��_ْ�ߨ�d$&��͕�P ���΃Q����~ɗ"�=ʔ�³��cʌ<E�-�UG >4�6r	.�͘�Gd�u_`K�y�BOgv�e-��Z�Rf꣰���?�~�8A��}ĴB�H.�i&Ӂ��XB���kV1���h�f�x䴱CI)���z�u&��0H�$0��y�p��Ʒ�Lp�#��y�K��T����-;}Q�	4P�=ky���q?���՘��j}oܕƛ�%��*��9l�n��fB���g����N����2T�0��U����"0%#����z���,,��C�Ŗ�~N�H�;���Db��$�V�R�Ǎ¼2$T9{Κz�D��g��6O���l�md�M�)n�2�*�O_L�2��3TtHI1�'���?nv�Lg^n��|�3�,�D����v�HzIwuO��j��٠V�	�)�Nc@�zQ���h
�k����f�e�Hn0�g��(�o����^h���+�n���i@�Z%�e���Ibpٍ���s�������!��L�Z�&r,��t��(*�Z�qăN���p�q$f���^g<���
��������ްP��Xi���=s1�2.����`c��2B'my!�/2*�t�p�sz���v�$��@a��~I�,�W��v�rs�3�kJ@�7���N6Ƨ��?��?�����/EfH�]��C��6��uϚ�S���)������6��Ņ�a^$�5Q�l?y�H]Zc�T%�q	)%���Z��b|c�E�}x�ϠR`P%��1��keқY��?!��`��Sܧ
�wF�okux��(&�)����J_�fc�<��z7dqh'�Igҡw`���6��hD:a+�f���f�U�c6Yf��ݹ#�8ر9�%.e�²C��X�h��rT���~�hk�FV�C�Y	���Y����6m��R�=��TA�F`,n��Zh7; �Pm" ��B���=*;L��*��}�2��Dj[�-��9����v��,�x�r"�hw���s��|���W��R��o���A� pB���Z}���cP�V�P �=�PN�W/y��jN#�ũWV�	�?��Aڣٍ�W���c��v}0(v�D瑞P�Ic4Ƭ��]�T��Q�"˲�����-��E�"K�/��E�+���ߗ虡�\³�zf��"�e�߿����5<FX���&K�n���20r <M�Ֆn>��2Ϧ�����C��%D6�_6$ǒ;k��_�&�?��\u�]��n�B�����u