XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k+P�\m'��)c�J��g.)F���CG"�x�h��>�G�A��\�Z֭�Z�{��YG�p-t0f��r�o���H��0�ُ둑Y_az��)�*���$�����1P�OM��-,z�1ⶦ��{��l��TR��?�ў�!����R��;��O2v�ϡ9L�����cВ��ĜW!(��Xȟn�o ��θ��9�x���8//��M�U@�44��H�ew��l:I�D��٘���ŭ�r�?��e���YX��5pe�C�~P��(�&�Wy���J�@�3����;(��Zn��Mq#%Ԡ�jx�P�r�Ƞ�]7�?3���=Ӓ���J�~�#�V8����#�9@^t$,[׈`��JC��=��|�G8+:aT�4�q������<WP94Q���-xT�ކ 97L�ȊR�O��T�(�X׍��w+��q(>����_a;م6�	JYFL�P�+^#�n6*��6�����+$	���Nh�k� �lד8E�
$�*�`����ü�a��<�����*���*Y#�}Z��B�o�k2P}H��l�
GȻ�V��L��Q�)K� ���B8z�w)��5��,�Y���)�c��b��A��?�l�f��s@�W���~?#�a��n(% t�����
~qm�+�pgJTk��P�/\������^�!$/������C���*��Ĺ[u�'���P [�H7y���2�d����CG��5�,��=Z�G�p�XlxVHYEB    17d8     890���)�	<�$?�/Ό����UZ��(���&F�(:�c��h��kI��!���SFiL2���Ӹ��yn�%�~7_T�")6�8�m"���x(��=��+�F�N����k`�B�+�3�1��pu���]�t?�w��Tӓ�?<)�;9�bN�|�E�kw�5��@�zWp����A�EG���|�o`>1)��PjgP�RbfEd{��>�
6rJ�6��s�1A��'JpY��gv�5l��QlkF]��!�/㕙��N�Mm�O���5���=7��[z�]��A2n6���LT��85�K�q���*����z�á��5J.�l�I�4o�w�2G��/ڌ:��[��>n�|��v�q:!�\�Iٓ`e�z72�PԚ
Kw�TV� � �)vD�� P�Y�J�����\E=�ǣ�aXr����|J�O��+il3v �dZ���+�j�FR�FD[0�VY���K�'y��I��ce�[�KM9(���F�>�i���zNe�������V�[Z%._V;�+6��S�A�����w`{���r�NK�pR����㪑NN��G���+,DW��ɂ�ko����u��(�
Ě(gƈ�1����|��� �>fTQ5
�]�6�Ln��ٷ��]�q1�.���T�aUZ�@�/��E�\���t���7H�ۏ�����I��ݟ1�2�3��2r�w!_�8�$$ǰ�}�i��4�C�Hӊ�����A�Q� �!}u礁I�!��+� e���O��/��d�o��Z���
=�Ɖ�*�Y�!}N#T(5���A�g�7^�)�����tWO��Xjqj�&œ��z�S8_���r����*:8w�Y��fD�4K]���q{<钋���B���xZ�([8Ң��F��#��o�/�5�\���=���_n��fV��Y�7�aJ��%��_7�@����-kz��:����,��hw{���P**M�Ń����h�%�#�� ��x�M�㑢[b	Kp2|��#��r�#�M(a�����)W03��ä��F��pjE�-��֧�-bHu���0#2{O.e����>����rض����B?!ߵk�����9�ɬE+)��<W$W�พh�j�k��H�Z���h|�`��e�ɩ�j��[�>�.�`�������4��I�|J�D��2��H2`*!����*���'����Xb㽂Aṛq3��{ƿg��;y?�c�Ѐ���uNgܟիBw�h�߳�[&�U�.�J�uAC�v�+��EPD/�
誟��x��+����Bi�
:�R>���$�g��.�n������������X���Q���$�~i�fG��dT(V�B{�/�kȓ�H��C���
PoW�y�1T��a��{�gNېe*��WD�D������?Q����o��/���r��V3�}0�\�Y������{�sl��+�p�z��A}��3^@��j�q�|���gB���HV��������c�L��������O�N��L�QZ����E���?�J���tD7<��LX�?q,�/����x�f�P��.��}ھ�����>����<H~T7��WF�����_��(o��q�,9#9�B�J=0��X;CP�J@Y�_{��-��Xޕ$����E�'�^�U�uĺDk���9��ȍ$�%�-ʻ����}�k����Bx�N��YCꓷ�.��|)��m�+w�f�E~3�U�%j����h��C�yD��8bp��?�־qn@)D(U�j����609��|JK��i����r���mr4����g��?QTl�����7�ʗ�M�bўj[�b-����+�dZ���l�����M�x$pWC�eh=cY�����G3ߚ�Y�Jk�˯��x��d��6K)�)�ɵ�ћІ��h&���U��k�!e��\��M@NQ�˩���*2i��p��?�z����p*�k���4�����>g��+6]6��pD����aSI晗�wc��k^Ó��O!I���MG��c�}�y�M��Ҫxԛ�����T����.+�G��˾���B�c�J[��Ҩm����Uܑ�f��t�2�8O��;����
%�F�y,��>� � ����q6�4�