XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W���\�G�C�/�D����A��F*��-$%LC�y5_2X��+�BN�d8�o�FJ�8�Ys�jJ\S��9#BX�w&x�nޥIb��2�ID� �H4�B�[�k������+[1g^��Uo� �0�[����`��읁p> �&�j������ �K��_��������O�ܿ�{Q|[�ϧ���[⮽���Zc�����2��!|f�s�ĭ����U�nr8�s%Kn\F��){�\7~(�,>�Ϻ�l-C_��_�1�8��	��3��62	fv�~���T���V4�k`�����ZbO�8�*������.w"�8���z��Si+�Ŏ�F#�����9�x�K����M#Y����g����2��V}��@~�ʧ��wɱ�����{%EaY�]B���;y~P0�K,şo��N�$�ۅ�%����6A�K ���j"*�R��c>v;�9����{�lV�DO����j΁��ݰρ�o�νۢC��3qox����l�K�}�W\����w!�9���u)$�QA#v�N!����L'-���Q��wA{���\&3���&8=w�ۋ�_���:��*y����L=n�e́Eԥ1�l�`�=QTj��mF��X�*�8��z�Z�!�J�=� �[����%�r)�XsH^�Ѿ>X|�R��L�u�N�ul��b��Fgq��H���Vd�4H �ͯ	np3�3lƛ(����B"����� '���#�[0^ҋ�ˢ�\��MCXlxVHYEB    af5c    1ad0�)G��[K�sZ�_�xQY�Y�&�B׀��p*�1SS/����n�E��D�.#�����^�͇��Ab�(#�yX�楹,�h���L߿����z��|^In�w��C��E������G~x��Y�^�#%xh��sɈ��]H�`�.�c�t(�W�/�d%1v�=�~�H��w�T=�"ہ(���D��Q<�^�	� ��a��3�Xqҫ췇���+g�2E����|F��u{�[����b�`�e�1���Yk]`�y�;ߑ+5��RT�\5܎���M�92i{,L��Lt
C�S��TM��|K�����Ϟ9�d��VY�;2%l�����4����Ҥ�祝j�s�I��Mh#o�ĥqdF��c�=GW&���S�M�8�<Lo���>����k�1�5��B0!B��}N���jk�(,�t�r&c�*�8�Cܲr�<�ʂ�T�(���s�ߺ���j/,}Xbz?d˄����X�Ò�� �-	���}�t�=U?��Wm��MJ9ꕇ$$���|�%�����" i{�c�ڎ7���.ƪ��`Z��	l�wU�� ��m�ﵲČ6ar��l��+X$�̕�EkͶ�3�&Q���6"{$�'�Z�q��������i����k�K�f���N�<WԠm)�!1>p�"��|+�֞�x��c��ϩ�$��j��F}O���G�]G"�W5�����ۖ����?�'I�2ʽ��}8�U9�� �Mef���O�Ma:��֐�.��a�ho��]D�S��� ���������`3�:����>���Ud�ϰi��\�{NZ��|���M/�{b|q��<;���Qr�?H�5�T�}��D�1�at����ۭB1	u�U���'��������tT)?�<��_!�b�~4��^曈ƞ�4��jzח��UK��9O+1�YD'���ިT�њ���Nٔ7��&CG�@��3O���h�=��ḋ2��s�sN�f×>*�8��)F���<�f�,�%'�,u���C<���p�t��L�D)Ո�߭í����ĺ�V�u���^�4��ŕਖ਼&"����N���5�?9r�g8�ݧU�y�jn��W�Pe]�Ȉ��o������j1p��R�<��5�VFk~cȮ��)���S�my܅\]�������l����6�J�swL�*���(�Ճ�	�po:�����4K�����pO)I}�D}��s�q=��k�'qa�����֯�!qp��S�OS��l���:¹��r�-a9S�g!�� �{���È@��I�)���Vz���s6)<z~�\(�3{[uK�+�a�GEY�����7�����o��ⱅJS�$I�^���?o�+���Ւ4�p��X�ݧo����s���56� <�5�1��Q���
3Ǖ�"�L3HR���naR�ͫrԐQ�D2�����n�QS#
�3ü4̛��[B*�����&��KHN�AKK<ʩ�D��Ű�;�.���aKà�8*A�(_��DV����1Ҏ����<x��мP��"��]����Iȏ:E�dmv�n�<wIyXnn<����./K��w��gn�|�bZ�zXR�d&0�,��J��ϒq�9\�)��Y�!^�&V ���4�L15�$0�߼��A�h�Iy5![~��5|��.8s��<��hg��"���̩��i2���kb��]��=��j�v�C��Q#^߇p��2�f�Ү���D��;�*���~�q.����fD��q��f�N��m��{8�r�=�e&�\G.�Pl��>�!�<Ѕy���ٓ���X0+SmƺE�F>T�:	�����e��,����"���>0�"�l���������v-w�Շ�~����z��g��Tn] �j\	2���=����;��Y��(����+ni��:��нVMuZ��ؽp��\D5��r&iԮ�X	�B�`B�'��D[�P?�ؕv�b���֞��3�Cv!�d�tG�\�xZ�pEI�\%�؆�-��2b0����k,�6�P��؆�H��G�����L�V
퐴�@Sr�{�S��L��, O�n�`{��;3�I�Z����1ѓ%H4p�I���� II����ȃN��Ñ�'	n�Q\t]�	�(Cn����� <HZ>52�d�;U~�O�
��zQ�t����χQ~�ĝy3�g��(��.��E��� �)}�����?C�l�G8ji�����G_���!96� �)B
}�q��H��<�v�u.1�kl��d���ʻ,�
�VV)"���W3x )�
�8�����Zo/
T̗��l���pT{f���իEC�������� @���FJ>�$A^�R:�r�������D�iT�B��{lꑄ����^u��7��4����J{�HP���]v�<ۚv!)�Wu��2��g|�ͦ�^%AY�	��h��$���|��`��X�	�ݾ�2I�� )8m{
"p'�e&�U�V���l�5����<@�D+Y1�yA��i�_PEb���;�L��EaK�@�]5īK/��F�eY��MSM;�,��� T�b<��?�:�Ⱥ�X���j�E2s�y��O|��=�7�-�6�+��Q8�=Q*�k��˂!3�3D��#גq�k�TRl��a��u��W�� @����=�؅�5����D�_�]�% [�u &ϫ���'�E[P8������N��W�a���Ysj���-AՔ�Jv�~�ǎ ���� �e�#-�t���k�twX���>�"�I����*��J�6�^���
��(�3��wlm�`c�3M�c��N������o�NX��.�HYwQ��s�=��W?.��a���q<���\��w�u�Vh�:��* ��;�^�x�8&��I����W8,z�0ET��*������=Q�H�q=���K��,ˇ�拓�_�W�6��-���4w|�қ�R����~?�Wd�������2���B0�[��AW���mz�c��x�넥v7Wط�@)��rZնI��d�ȟ�in���n�N2����ڬ�,����22^�=���?���܋@�P�T��>XĜ��l���Q���0� D"��+H�-T-w�s�C��NRpư��(K��)�2b�{UNJ�E�u�k��bg�vlRP�z@�Fah��!b��F�o�q��O��$�g=垹Ŀ��vņ����1N���3�Z7�y�>��,\��ȋ��Z��&�:�i'��B5��������Bt���n@z��7�J�%��q@�kIi��CAV�L�/�.HR�Mo_σ�~���'�LR%� 62���mO��2�k@�i�V��8M���'1g�k�H<EP\fa�Q�C�5�(�]p����6b��|�P���{M�������1x4S.c[��Q�d�g�b�����~��ԉ5����le~){ڋFw*iR����*��F}[$�U�5�*�`怒ؽli��HZ�ӳtgn�.���:f�l��w�MN���ÞH^MjRwN�T���ق:�[s���J���w���sO{�{� V�!=�4���x�~��t�#��G{�E�LY�d@?��S�*��q��<n�ع����;�&�� f����j����(��՜S��I��e�5�Q\r��)e��ϡ�|u:�hݖ�k�g��]@Y`pk�
�
�<��WaWb;r0gq�l��*m��<t����jedb�K�H#��*Եh�^��ߝ��Y��H���Eޒ-�s����w���CMx� ��.4��wP��ܪ9�: �D;c�e�ơr���#�8��lzO�m�g�m�ޚŋ (���Y��.ڢ�iB	V鼞�ҍ������(���������eZUƃ�/�e]8a��?��:%s7���X����Z���W�(���aw�~NK��)�?�'�;O�!�I�]��(q7�tIshV'[ǌ't׽�h���E'�,M,1ٸ�����B뛐�RDod�4����1�9�Z������rIJ�l��TjC'$��W����2����-ޕ-�-��jÖ�,�:��X���̼^zNy�'��k&����x�L��E���ddP�Q��m��	 ���=_mr��b�W@����T���;���ޘs���/L�D?��Z�p�Q��X�S��Y�h�XpZ6�9K��v.e�����dW{jaz��O�RC�}�Wl��d�>�	.(��b4N�8���q}���
p��B[�ymX��-�=AKpIyZЖ1��B�,����,,f�?D���̷Yݺ̺���q ����\_�~!��Ñ�2�q'#�oa=�)x�h��K��8����3Tmt,�9��;�3�Y��-}c����4�	����o�Bu����SU�������D󰄗��슇J��H�Z���#�	�y��6?̡�{TGZw~d�Y��փ9S4��[�	�t�>���l=<�����gg�z���r��2H�t�=���jR�hvL��jNn� v���S$��e��5X��syK��<�"S9�%4�ѧ�7���>(�W��y��j�Ş�HFhi^8�%����x�T� (s��ng�g*2�p�|5�,M�r0>MB�@�*u��^D�L0�E�N�� r�=��|R$*z��'�����%p��/$��B�UR���Hjڜ��I����Jy�Q~$����A���\�4M	����c�Unt R�7�`�+�r�`�xϫ�u�wyρZ���p��UZ�74pv�~�s�����-��nQi.��ն��qQíE+�$�\*��>T��������|�oi�(��,`�o�>:��j.�?�%ZU��� W��+n�"N��"P����&@�����9Ȫ*�w6�;m�.��E]�b��kV��nt^i�"�d��<�LD�t���*^��˖��;�R���k���b?'N%�@=%�N*:�r��U����I����b(lRz@�
����O�ÅXh�=�p �j�os�<=�e]QX�m�BCCʯ�D�H188�.jFł-iʜ���o�2si?���r��:!\$( ��*4�q�.�`�6�^�d�}�������O����xD����M��ſ>l��g��@��D�4Cl��P�)��[#@X��v�v��/�0v`�(L#�0HO#�r��T�OB���aF�+mF�e�G.s<�w�Ό���t���2c���<7���u���;��`�j�Ǒ�)*�&iػk�0 BS�<�-�Bh�M+B��	�L3�S�k�&9��4LeV�!T@q=	WY����c|g�������A�H�G��1�;/|�*�dNCĒjKt랓�@뛭%�����ӓ���o������H�{�:!Y5���,�6����0
�ծ���%t��=��;v�(y���+cz9��7M�����HI��2��,+}���4��aK4�Ư�>�&:-����Hݨ=�ݪܒ5�}�DM[S�:OL� �N3^����C2���R=ʔ��K��D��b��Pۺ9�-�3�~>:�zS�K���3��1g�yﯩ5���J�ثb#)��j�Qk��!�3u�X�4^3�d�x�/��(������] ���绳��+#(�C�� �u|�W����qx��e����D���K3wS����mN������|Bm�?z>���}5�i��q�O+~�"-���آ<�<zg�4��4��<ٕ��?��j;����+�s������`+]�2�j��͠���Y��Ч�d��&jBR=�W�L��b/� ګT��PK��}�ha@h�&Q1��+͚���hf�]
C{��gM�E�b\ �{?"9fױ�u��S�Ix��������3v���Fް�a��J���U��ŴW@����Ą�y�	�J�Ur2j`4+p2H��p�ҕ��E[ȁ.��!�&�n빸�hyR���P�
C��q~68���p��Mϱ���Ï�Jl�����Fs��:��U!��Ʌ
�X}��9xy�L"��x�AxK���ǡ�u�$X1.��O��1^�~�= i�n����0��_��L�����D�D�6͑�hj�����o����A���gұ���ЄT��O�3_�cV��O��B'd`�}��l$�.����~����!�q�����Uڡ|��+ *(����V��[dw56=u�i�l� �۶g����l����̞�:�ؖK�b����ۀ`o�k��+BД@D Y'b��^[��w+�����U�^���2�'����#B�j�Ey��B�W`�CO��*GOq~�(�^7�"Ҍ��|t<~&���S�g���=nu(��̯�/T	 �ď�"�s�e���Y�Q�Bs�z�C~7| wT�_r�|8Fȓ�Jbgf&�x$��Gmb�|�.0J�n�s�v/����F9�e�r���a%��w�]�L����T�j�0eT(?�l0�,� �呶%�Ů��PqTC�BۀD�o,ӧ�[%e@�36����g0��O�tEzQ��� p0s�A@��z�Dg�As�4�jfت
O�(�ڨ�L01�K���5\qW2#�kf#�}̧��aiyŲ��l 6�%�ܐb�%�)hdN�<i��D����2sYF��D�|����X$�m�G�T�c�(A��"��a��[�8��c�"�8����,�<��"�1ǘ�Ѥ{���oG/.�Ǳ���Uv�*(��,C������� ������b	e�5�Q�H07�;̭�Bh6Lص�5a)Ķ�A/.�?��_�Oe��ht�<r�ڸ�7��}"�^�����C�n�