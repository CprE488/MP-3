XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����7�W�({���bL��7�wO;+B�5c���ԙeN��,�����k^%)&�ڐ̦�'n�&w�Ii3ޞ]\�Aw4F�T��*�v�8�F�:��$d�WT��j8O�/G����u��;Q����5��s����Z����#k쯡�RF�b[��*�2m˿#�*����k�޶C�3����K����G�Aˆ�DްZ����`@:����w�,N�o.�^�Mĥ�B ��sE��р��
#�3ĦIS�����'ow@]*���ȁwr<�9d��w�ϥese�H��V��soO�J<��`s~�	9������@�򰴊6z�Ż ��s�=,��;W�t��Yzm�-�Qn����E\X�W�H�IF��{I�v������`��U&3 (TQ>�'��h?�I����-�)���媡d��YȐ��#�YJ�gP_¨����[�F^t�_|�6���>��t�2W^�-�x����r���I�=�i����kkx%�KΤ%�*���Ň�J��]�$<�8�|3l�N*�����ʄ���e�;Z�|��-ek��)���(�tJ����j'�������V����|�ı��:���6�XЃ:9��+��Wq�|p&�`x.,���+�	����Ë5�Ħ)��jN���s�p��zY��PS�O���\���G1�#����B$o�>��8@�����ɽ���K��Qsl��~����,8�U+����XlxVHYEB    5fea    1830����!%�����z������]��"+L)@�L���
$�����5"��c���U�<}��D�+��n�� 6pf]���
z ��)Qųz��q�Jܾ�ϳ�B����^��!����x�]��>�������H�l�
L�(r�m�ՙ��w��&/W�i� ��0��sJ�G/6(\N��p�@����QZdmH`��7�b�h9H�&����T\u�Y9�|�9��c�G�� ��u�;(�fEǾ���o3鏴�����}��9z$C��W�x�Թ����d";x��]���*)!�&��V���Ys�2�J��g�f[�8S�c�)��KL2c2�Q���[��$�x=j�]ԭ�3�õ^Vrɓu����ibR��H��!� Y�imeⰘ���T47��˞��y�xo���B�7h��0������;��0��6����՞�N @W�M��4�P^yE����Bq|�́u��a�ړ�7p=�P�1��R��gQb�wf/f�=4�?�WW24(3�\���h?��-o�Eᷛ�h��}R#��冇
�)w��lr2i�@6J,���^qM=O�%�y�J�$��	���vc��s<�����o��6�|���$!"�"��D?N��w�܃�MϜ� .
�6�2!	B�մXn�P��cW�E�cK���c�K,N����"��*��=�q*~M�IV�PnxX���d�T�:�h��&FttQ�A��N]�E��~���ݠ�ѿE��FUȺ'z%R}3�ӊ8�-7]@��G$�5���Mp���b¡��xu��r�O���}@]]�K�i�P&�A�������R���q�}c���ۆ�)�]�gB���f�7��Ȳ2�Fjz�U��Z���Z��n�{L�����ѡ���I�?D������Ke߭W������ K'
lQ���t��H'J��=<�T�5�	�8X��o��R`��-nǻ(��� 7l��I㝥O��_Հ�7�ʛ�D>3&d�L�P��0�w���^-�=�Y���w��\.]��9ra	è>�XhNO�(eK��헤����OY��y6�^)�CT`��(X�oݢ�xԵ��ɼ�eP4%~]3iۀF��ʍ_B�,�,��}�gi�B&E����6�˟.�1T�ƉP������˓�h��Û:_p0�(F�'un��"��py	ʪO��j[��=S�(��U������Gs�yÆ����mA�Ʋ-�!���b3�+�~}�`�h&�,K7|�J������ u.��BG��m�zH*�\5w�����56�b�U���?2r���!�˅��p�2�0�Q��J�&���L1�
�d<B���~�{���?}�\���-�������FZ$:e|��0�����k�l�k��n�AZ�H(�.����2�>!:v��ep���x}���~%�8<wP�ę�~��,5܊O!z�U������`j�aѦ�"M.����_Ђ�&b������;�(ڤ�yr-�M�蛂��'ڮ(�/qn�\p�#5z'�ɼJ�Ϙ�U�l�0ůi5A���J��ߑ�U���دX�ڦ���|J����D]�W�N����T�J<���9�9��&�B:~Aa����+I�Z��~�R��5Q 8_��0�!���/�U�L*3.RMB��a��T�$�:�Y�"�r�u�%�l8ql����%��h&۾�|1,�|����v+=��)����}RD	
����ɏ\� ���t��޵۸)P������y6�Ɔ�eg;�ӼZ����}A�~�����e �o<�[nl���)�.5��+�{K����S�(���V~�Rh)�M>��q��N���V�.�4�R�r�t6�FD�2$��4Ɂbڟ2l��h�A��%�Z&����ݠ�hkA!M*s���BO�2S1�Jߩ�A��IÒ�c�]���ŉ�ڬT6�r�����ҥDiU�4˫4�(KOc$�^n�7@g�s�Ή�k�R��$��Β��:;3B)XG� ŝɟ�m�xG�?W��%����4����_#H��wI^��x�����6d^�{��0��Y%��#��}�M�c�d�ʲ��� q�֕�LQ�o��ĬL|��g��xJj�|��2ǔ#:��w�Tol���$�~0qb,��|�O��?��������@�&#�5�$���@{'m��9�M�y���B*ji���l1
m��@js�G�Ce���Y����q��'��l ��8���=ߠ�
��J��6�aWD&�A��}�7������g)��{�!�H�
��5��)g%!��)��Յ��JL#/�7�?�rj�Ϯg�,��eU2UcP�S(��/֑��t�=���7"q������DҺ�jp\�>61s34��1�������}� ��ED��S����6���W��p�f�g�(�ӯXY[���d�_ ���"�U�G9Ve�vU�Tq��BC���Tc8
�r��/�R��ޑ��x������q���׭z�G�<"N���`��ʍ�%k�v�A����;�m��m��bN����m��9����G�w��8I�M6E�.s����7�{V�����{���h��<�%o�;�^6Hk��K���㙀�	;�$uhl�n��P%o�$��69Ҹ��a0�^ܰ���)���6Le hJ֘��`N�:���o4�?���X萆�X��ƴl
�����1;��&%=��,m7�zn���4D߅��$� �������l���>Z4�:�K��7:a+E�E�ص�X
i ����a�����F|n' ��RQu�$�n�Ŕ�R>�VsE�X*a��>������2��X2F�d��jI�0ד�R�DW����
{�.�!C��w��i������.Q����zD�F� #^�:EDUb����E9θ�q���f���8�6A$/?�.��)�t 53���4f�;�a�U>��5��fº ��1C4���ݿ�����Ʉ��*�`��%[�I��%���!Ę:�b{����&�𐪏JՔ ۈ[������t >m��v���/��E��}�����g�0��|�΂=�*�k�.T$��!_�,;_��E�=�z��j�4;�EO� ,��G+s�Hu9䤮��PA����30S�@��>]s��5�<ø�
�C\���R���xd"�f�t(xy����ijS�(Ἦ��`߭������B ����d��&��%	G�sucU[���$�0�����_�Ļ:)�����t���;��\�?/��gTSm�9nܐ����ȾZ�~5+��H�'N=^��ͽ�ji��@��$����̪��'�~����b0Ј����%6vd�p@nKÄ6bm~��\���>�)d�^�л��Je��0/�I��4�k�ތ�j�����e����ODG0���C��L���$���%@_N���|��Ҋ��G���x*�l�R�V��5Y���{��2��YJ�<鬮��5UF�s�/�n���c�Ъ��&1�!ҿ��c�в�j�!=㕈[�"�hr2����`�)r��2��%sZ��l��}g��S-��~�;#��0���if x��ܢ�f�����r�@��!�w C/�8qmw�
��,�1/�znQ���e2!���ѝ����(��s�d��^q�mwzDoE�E�Q�s�:@{�L��/��u�mr���C$~��8��!�$rF�9_;���$���.�s�˱w����]W@�`��II�ԢJn���3���zv�4�l]�Ǐ��f���e�ð�p,��O9 a�Y���>�,wڰ���oծ�=A���xw��u���'wR��
;�$�K��7�rៃD	�{���gx`'ٵJ ��ȃ�K��9��&ʤ�2�q�6��l#~��,���4��]B\Q�.�����Ce*���-�^���;��W�Q���O,<F�rċ!s�m�����/EO�5wW.c�V�F�����e��Ԅ�s~%��d|�i���դ���.5�6�l�9~6�Oj�U�~���ozp�g��/gp�u4��k�ؖ�^5�Z�IC�l����$1���[��+�H,���jIN�s��R@t���H���H@\g��S�}�+��<pb�j=��ߵr=DS#T���q�:�i
]���׳ݫ���a�glٖ��������#��"��&X?�Bc����Q0�tk`��cX���F@赞.�El�}�l��/_K�Hw�0<%�f)�_M&^���d8=:����c��D/���c���V��� N��4}���⢉�Wv=�ȉ�=�l��U�]Y�K���>2ݗ��RuM�'�mp�*���Je,t��:����?��1X��������}I�wRa]zHM��#�z��%Ks湑��~"��O�Sˉ�)e|�$X�!���U ���T�Q]��g�rX,E[����j�o
�N�BR�D�%P�\זhMi3uz�����LL�fKv�U��p,:b�p��U*u��_a�,v>VP
�j���t/5Q���jԸ�v� Y�z�
��\E��:X�l�48��H+��.�z+����w���Y�Ħ٩���<G "��%�5���������1����Q�@A��XE���0- Qy���8�q�������z=Ѷ�t��qW�z�q�})6R��H��W�p��[�d��p,����$���A�b�U���/շү�b(�?xe�j��)�S*N���ӻ�H\B��ŶdX��o�� �R^��WT��
���wm��$ׇ�]�1��i ��l�]G6�~�� :|��/{Z3��rL�
U�d�J�ڦ��{,0����zN�
�)[�nC 8<��H}?R~6�D�zK�MǕ�>��ˈ1�s0��W*�u���v`M��l��|z�=��r|����v�=e���W+���bE��=glS�=m���!�_��-�ɀ����*��y����9�mwE7A�oUB^���k�q"n��f�+<�<w]ݖ,kq��#��+��4S�M��A�	_:cn	�u?n�'u����H�v������8�c����Ѧ�rb�|��7����;-/e��A ��2�U��YÌ��~���F��]�.�ί~����4r	Ԋf�ټ� �\9��<I��>�	�P�N Z���$:O�O������qL�ө����a&G��_�`t��|��lW6b�oKl�_@CY�N���!A�^��C%b�($7O����%�s�u���G�&�ZcB0�����i��I��;��ܹ�7v��W���,�Kc���z�Ŀ_͆�랬���|�H�u�^oMp)5o��{�?k�E��E#�����JjTVK��)���_sqj[X�2P���J�NC}����	���L��0�NPcC�޾����������,历8#fۖ{��bP��9�*nH�VF�)�OcR9�hUq_���q갏[/��*�N�"ؕM1���āM0��p�ba����^�����������Z�<��r��z�M�&+��Q�O(��p�*7)}��)0&�U�$W$Jŭ��=O:M1�b�~$����cT���L����R�h9�3�|�ٱ0�������uțϚ:+�	+�9췩�s�i��8*L'���{�����!�ڔ��[8��y�s�C �1j.�?Ǝ�d������.(J�j�I	�f�"���db�?�NL,�j��0�����]����j K޶�%��`��<�I5�������v�"'�L�����aWMz/J�.� �C�����$bW�wGU��u�UKv?Uc���y�V��E.��E�仾�z�u�()���nu���,��;*����P�,�����ۓ^Q*FyK����,ѼA��M%"��'j�8����4�W���IF=ӖP�z�mGߞF�{b�[���W������a���'X�4����O�a���̿�����iη�זi��Ԁ6;�A>f���1�l��GO�ɱW���u��&�U�� ����r���[�����ye+2���#�����w����hA ���=�k�w�+�*J~/:)�X�-�.���<J�ʁ
����,�I`�