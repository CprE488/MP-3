XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������Jap�"l��Ѯ�l?�p�+a�.-�}��bI.�HZ�"�O���|E��[����p��Q�p��5�!U7�|m0����#,P�M8�W�}���=Ğ��g�7��#�u8�
P�x�"!$ܭ}�ʄS9�l3�̵�0�z����4��)����@��o7�UoE��!N���l���A$R�p��:;y�{�X�w�pA��ײثG�jE�k���0'�������1�6�&����<V��v%�!���JH ������BEt�6�AhӸ+�y!�J�*w=���UF�o��֦9`�[vX_���RH�X���q��+�ur0o3�U�v�j-~4Ҩ�W����7u�A���1hS�3�.�G��
�AX�-�Eɐ��|x����p��W(�z��;��⳷����.|�GtrA�vE�-b/���;����`�O.;����ź����,2�4:��z5����EȲ!���K>��s~� ��I�K�������)/�� ��,}z�Q�="�~���	TS�ǣX-w���@m�aW}��+.C_������h�&��!f�wJu'GA��͑�e�]Gҧ��]�@�����������L���F�*�2�%�: .Kt�:iNr���D�Vk��0�)L�m�ѳ����u��Y��V�	�=37Q��R��{�@-Ʌ���~���豝s]���:�C��%`� ��������ЀA���gYi#�&Պ�8s^��]��&D%34/XlxVHYEB    b087    2540x�@�W@RQ�Q�eK�M��iȔ �\A�K��?d�6�p�H��v�(������P�Rت��ɒ�~��bE�mij��H4���,{	�+P��*���yݷ�	�y#�x�#j-��h�r?Td���2������9������Z乙`ֽ�$H82��*��.�e�s�9z?�Եݸ�iw����ũ�
�ݯ�V���[�Ԡ.ui�h;���k
*�4���=�=;��"�dh�'"8�mn��|R��⑝�X${���w}����[㐉p��{y�"K�b��q�����-d2b�]�wά�t�Y��� �˩f쯿�{�N���/�4Y\	.E�O�D��K/��v�w���%'�4[�ɍ���ɥM�Qn�[t�u�O&�>����QP�x��lN�1�U7�;:8��z����k(����ʢ}e��x�ے���(_�fE�� �[�����	�dN�̭�gމ"���l�Tɖ��k����?�o����sm�H_˥f:j���<I�'�N��0���?UYޕ3 �b;6���!�L������ȸ�z�j��A��	�����4S̕�{CB�=��Xqّs����2�Ev4ۂ27NQ%�go���LZ��)���7~���j��'��I'K��J�X|6%�{��L!�{ ��SA�������D�n	��b���Қ*+C�Q
b���|�T#�� �֘�����`1&�Z�jIqc�a�#��@?Y��������?Bn���n�<�
"�¶�l֍Ļ�H����fOo�"_c��/�V:�:ab��wf�>�D�(¸P����"��>�O�z.|Nsx�Q��@"U�N������s�_��/�ʔ��	��C���3������6���1���q#��NY�{����)_�&iS�9��뱺
[a뚡�r���dB��p��bވ�9ϲ���X
�0_V���=Z�ޒ<�Rw��9��~R�M�͗�G��,z>��PaF����g�Ϯ=a?D���̨�V�tXϪ(뤩5zq���|�\�!��Т�3nueQ�uȧ��cF��
��/Bz�d����c�)�s��Y��5;�s��P�84GZ�cG
��=E}�M�|N�瀨��v���J�����N&qǼ��ZCf�5/)� 
H���q����;�^���O��ů}^�~���o�K����H3$���.b������~�ɖ@Y��>d�#�W.�R4f��/�T�Qy��ۚS� ���f����9����V��j��F٘a�<�<�-{"�&j���'�ZC��hH���X  :j��sƸ,܇��+�5�C�Hʰ���ny�aH�\��O��dm�4�wU�o���pm���qA��q>�}��|�K���`�'�/��~��x���A.9�7�?��d�!���C�PvaB��ި��s��C�	s�j�o�k�����;�B��]���F1�U�L�F���_	 4)|�+�DI��9y9���M��'#[���ֵs/Aܬ�ʜ��&�jN�*S,0D�a%��c���XH�Oُ�P.�D	��]r2�k�89�NL�� 
�2b��+>����bL�T35M7-2����r(�Rӻt��\<e�	R�֑�R�]F5%µ�1S���3�p�����$K1�s
X��N��0B'8r���eO�J��v�Viƙ�Ǆ��G� ���r�鏞�k�'#�߃��X}��1A�̙7������t2��ג�q�r�xg�y1��&�A[�n R'����l~Avؠ��r�G�OƵ�5b���*�Hʹ��,<P�,E:��c�/ G'3�v�&R~��艁Ƕz ���\b����K�	��8l�)!9p�I���9b���\ |�8�^�	���u� �0k�6(\�^&�8�R�s�� ��b5��,$���88w�ra��yJ%)\}��_����~���c�W���F
�ȍ�
s΂\���kڬ�s^�0�@�@��Ǘ5�V�q����r���p6� `x��1t�?m5M�JTN6,�l��K����܁d@��a�K����m�j/k��D��/��RVPNu�j���4�$k�䣧�<~3A�M�μ;��j��
�0D�+�aX�=L�yC�3���GK�(��p�$�0p��3ܾ�� 6�C��#����|�l�&�����w�?c��iEJ�ez�^�9֖��Я�DD��D��%��H�I�T*�"��g?3/}�:���Ó���
)�Hd������|`gR����>��E�u�bZ�*�Q��@��5O��X�������LdG�6���[p*?�*K�4�U]j�O�D&��[u&&�]gE T�% ����x��-N?y��q$a���Xl%ҹy���XW�re�����q��V08�1���e0q1GNؿY��d��j���;v��d)�M��sG, ��S��D����NTӠ���z���T�,�΀}�Ɯ	,Z�rKy�&����lW�E�Gl
u+~BR�7����ӬS�=�s�N弆�vn�Y{�ԍ��=��4�np�/�)�UѸ6�?Å�y�Sm�Bݴ��׎{�MT)(���Z�f�6�/�k^����G�iǉ��� ?�Cu�`Y��^�$|�i(�$����ˆ���,F�ᐉ����g��8���1F�PWf�L{�Dw!g�J�b3Pg��sYn̅%����3�v���9w\��6o�|�]M� ��i�w��x�&#��6��L&�Z�s� u�6���3��n:�S�����X�I�R��j�	,-
�7c���6�"�i#Q�hԏ��MQ����v���?Мg�h�e�S�5��h=Hm,e��\��i�r {�o�g�%iՀ�����0t�R�l+>��JI8�p&�3�nFN�%
�$�YҦ?
I�Q�(e�8ߞ�������%
�g k�өw<c�T��N���!Hy(�R�Omy����05:����\���S����v<gkka��_$T�����n�k���3� *��mf�:)��js��.���G�Q�à���r3��<��C$ g�9�aӶ�)j+�7rn5OB�[�4M�^���o�E�_���#�Y�6M���%��k	�kc�<S��t�0KLm1.�+�.�#�)���$�;�	6�&xx7���sT0ٕ����!�7Ѯ�٣�WvN���5�8�+fM����OzR��܃���������sY�܍2=^����B�ӎ��6��R��km�|�:�l�7�nD,�	�F)���x�k$�mL��@�%O�{T��tc��)*�ٲ���O���)�q8\�mػo���r�#�%3���Nh������[Q� {�T$v��m��j��D��%⧗O`����}��4�m�7Lnf`�(�]
�T)���Q��h�Z����Ҡ�����L�݂��%"���w��a���d�n���6�����Pf�`�/	�^��Mj��6\���p^�n=g�A�d/Dz1�Ud�O+'
�!�	��z�F /l�f�5���O�x�o�V��|�B{C��ե AV�8N��bfrY�^Q��<�5���e�l�ŭ�W�7L��~�%�H����^EbR��}|�ky1C�f�[�[�2�U�i�3�Vǲ����.Y�!J�K,3f�Е>���B+ZQ���*8-�B���Qp�Z���R���`�$Ө����z�"��xZ�#Sb�8�E��N���?��p��^
6uaU1�f)�b����kO/��Qm)���p����$,|������_z{�@����R7[qLȫ%X���;�V^J�#���5mH�޳o>Z?���{�km�BR�N��h�m����7��	�M秏Z��	f��5��@F�S��A��fq����y�;'����K{�O�	���6�@9�*��
b��Ck�;zuhw!�Bm��rgbx&�4�_��k���:���_`��FJ��Ă[���/�]J�hֈ:�
�o,�aj�el��s����#R�T�R�sd��ӆ`���S!_��G�x �ы�k=�d��8��!?��]��y=M�F绅@C��P)���#\�6{�n�l?��g�I|�~H��HR��~�����g�x������7�1�޶�0��8)(mj򧙹uS�Px"��D��7�M��l�Q:tش��NG���;�m�D0L�x�׍'H:;cPkT�[3Zu�-G�	�йQ�>�Ϡ�;��^��@6�+���HK�����$����dWՆ�<i�����1�8M$z���X'{ڕ~5LA3-:�K�8�&��_\��K׈�4[��_�Qw9��C�W�,��� �R�d�/�@�5w����B�������3�t��F��̰�s>�)"�F+�<zp׿0l��bl���5��`D���!���3��&��dS�A��}"�0���"H���r>UGٰ&��,�gi��U���K��n�r]��G�ٖ��5fn@>)���
�`�KP����+�R�z[����|�q��O�-���v���O蝨���pYKLDTlC>�JV�u��Åu�����G���
����2R��'ج�����l�D�t7&�s���smM�C왺�<Uj�;�UT�_�QT6�
�B���vsu�69Mt[��<*$T�w�r�A�T�';3 ���4��I�]���
�d$�D����`aq���kKy�wa)M��:�G��}�٨a%�3��H�`=-*"�#�w���T�A@�h6!{6k����i$��*�-������1�o����󊹽�S��S?�S{�Q��fע�<?���9a<T������~jh�塊Wlp׊��fOz�WeSm��Ҿ�?�E0D�����-��O1@ι�r6�>R9}�x�ic͕��:����Ѓ��t�[���E�~�Q�~`qۤk�?����&ĸ��`��b5V����뇳�TLt���	��d.��TK|�h������֟y���|[J�����!��ev�h�����J��%bz�ӫY��u���S��~��ar�JG:��8�E���L~��)f)O��Ǵ<*�^��l�]@ћD"@iA�9�v�	�ɼG3I/
s�>�|�ߟC\W�ף��;a>�������Npn�$y(�˴����s�d�-���M�=�7�4�s�=K�7�%GF�ˆ�L͹��Vm�[ig�ۣ����X����/�%��~�M�
:�vL�7*+�U>oG��J%Œ��i�=����
��vR��D�ϛo�N't�����B�9��=����#��X�SN���[��h��ư�Y��i�k�b�v���a'��)���O�2�n��?�ajr���t+}�d�����=w�����T�_���^��,�g������:�Dڪ&x�=^���E���2�)�F���1����i���OGL�^�PN���Өt��gP��@d��C=�ti}��<ȹ�(H�t�X���� �*��'p�TI�3����E�>Z���Õ%����@.��$O혜�����;ց�hy�*��\�{p�2h
�x.=x:vyA�/={f&�$tη��e��j��3	�5�V�$Z�3�Y������O�U�e��z2��"�C��CZ�D9��fy�qb�4��c//2��k$ۮ��LR��D�k8<璩S��[��F�D"Nƛ���8�#��e)H) ?y]�����p�HtT�Ҕ�J�~��bv�%�>���)���]�];��&�A�;�*ř�;I4�#Tj"
9ʠEA��:KwEu-tsشf��l2\KNVW�m�M���s�����e�^O�«0	���Å|3���8^ ���0vl�U-��r���@�0�nPdBF�~� �>�G�j�4B->�K��J3Һ|R��:s�i��s�P�#.��+�)7.�QR��89F�������A�����?+m��s�c������MZ]e�����+�96�`Ǳ*F�gb�Slǅ#q� �w.�e�I��N�tji�k�~����X`泜M��jK�u� �-�jϷS������%Z�\�s���� �2�8D�3�0\r�Sc��_�]NdR�#�9&��p[DCT����l4�N�JF�S���ݻ&��������27�ML�ʚ����F
���>�%4���ʿ����@�:��'�e��)u��:��{��N+��o�`�kUZ�$b��
���~Ī��.��M5Y.���΅��r�5]�Wi���d����7v��b����t�9�s��dhNJ�0��3f	}1M��E� 拓��N�z`��ԉjz=XS~ �rf{ݑu���9���4���Od%��9-h�;���Xܖk`Rm�\nb�%7i��YJ�����V�FP�d�RW�ȎΘ�ja��3(���=j(�B���S��y"�{�}=���§	"^�&8�:���	�ݛC�iЁ�� Ax�ƞ�+7�z�isF��J�H~�u�)[AB]��+fY"l}I�����LX#ެ��ys�IL�ǡ�%�r
y)�~��ӧ� ��!���LٸC��(�m��O�y�A�<�JǬ7P�*�T(S��8��,�fC0����V�Z��\'hܑH"��^b�CR}�A��(Zz���+BǄ��E�="�L�V��v����"�4��TǹZK~G��*x�k�X ��>�P����p��L:E�u_!��~֚����]8v4�<��?'tY���c`K�Irf�c�{k$�ǃr	��P;�=���D�X�u�wG��]��	J�"��= ����Ip����5ؓh}D@C�C�Q���ξZۗk�� 5V5�""ǹڀԷ�06U1�����˧���l���_��j�[6��炲� �nɇg�*�9�^vK�����*Н�I�y}󺳒���"H"(5模�E�vc�{<ᣰH��ڳ�cS�HU�l�fa�R�t�LnR�V%��M��?�vc�k��؝�;����Y��G��,�pe��9?=:#��~ޡƗ��&b�j4�,���*���@Iu�[2
J#r�I��Dh6�����w�HѠ�Ͷ��W:U�<���į-V�oNZn�%���=���}[A��'g�^�Ђ\�����*a�.�����K%"V�ٟ�X�Q؆�yS=�"s��:����P.�i�`���.ax&r@��^�J����3�{��}2|T�Y�b������iz��ӥ�jž���}�j�k��{#���t�]c뱠��w�I,��=�X�<���D�;���Q�4��S�c�Z���?���L�;����R����L����O�x��YD88FQ	��~$[Z芊2쵺����㙱�G�gO����L�k����:�xJ�u�(C��X���4�Z�7�2�EH��%�Q���(��*��w�"bf�Q�G-7���bR�WDzw���KŒީ��c!��k �^FHZU�x�o*;m[��6�������-�N7�[%L�_ ���̛{R��n�E?���y��s1^|*
Q���&��ߍ���vQ�F����'�tki�W�T�X��971'�Ѐ�etE�TS�%�Ps���dPt���<��ݢ&�\��}����Qp�R�����9��e�VI ���D(2w	f�F���񼧦����0�����ؿ��b�����Ya�ʩ(9cJ
�i�<��m��lb��I��
w���^�Ia���I�R1��`�*��?��I�I�,�p�_�k�{7�B�[�i�+ȓ�7g���2�GpC���Tm�g���<�V�U�h�Q�ڭ��2����钾a��#z��<�u_=�}X��`-|cG�[�����⃒��t�RM�j4��T��	D����k�C�X�3�,z�\?G@	hu��Z�Њ4��*%�*�	�<�o�����OWZVOq�\[�:7� �I��� \�_��=<ן����0������ѴK�@cE�G�Y������ͨ�a��@���ᓳ�7���N�(�	��"��zMqK�Ъ�|�c-U����WR�IBK��%��W;�]Q�Z� |�~��U�ӯ��F���eB���Z�$��Y&��u~��=Y�`=��w��a)&�,��.��BN���K��,M���y_�]�*�&��@�9�%�w=k%2�Gc��y1����WAv���\/˼Fm�1��af�'5#$Sa�*x�jW��"�bt�[�|4Gha�#  ��u���D6�	U�Y�Ty͌�;ݗ�T����`�O��0�~��i�����y�?��QyYG�;��M�@m�� &`G97��g ^L/`�!�{��l8�/���>�o4%�R_aV�Dޥ���?jtI�e�sz�M�,��5]�b7���5vraB����h���F�ZT8O�H�w�|�0�Uf���&��)n[جW"E&��D؊h�8���>�=ݖ��(^�^~\���t�����7�0#���jJ�\�כ��v�4]읿R��I���o�����庉�e"+�h��1�~�
�A��Ź��V�r�y���	���j��v&}�)��H�J�E>{��o!5����2-f�a�}��Md��42��wi^.˻���{&a�j]�<HwX��<T0��(y�4-���e����g����A���9#@��6gZu�'c,�>�=Zɳ�g�x�{c���
�:���]ј��g��T4�7*�5Zl�c37�"lH�9M���ʥ�D8�����_�����)0@�@݉9ގ������taJ;i	O@6��꯱#�U���j�����XW��{�+���9�L<Ę��h.fU���ڤ�;��P�e4lX�<|*N������Dڲ�ʬ^�e�"N����R=����r����1�$X��i}=���Wi���ҵk��S�1���O������Mt|wǚ����?���w�����\�*/�6�mX*֤<���8ßt����G:K��ْA29R\��z ����1��ǁ��d)���ð������ ����Ӊf8�۳ls�1�#`�XZU��W)>�:��`�ތ�4͆��aw��4�YK��{h �;��F�V��M%=b�ZqbyiL$%�5E㘉o�^i�Sfs�Y4�����]�]79:�3g�D��|o4\�eV4O�1�����-��}�AU_��=o���.-&��\�xtȆR���iK�G�W��\I�Ҁˑ��%�W�᜚�d��=���π{�DN�E��N��	rϵ ꬗_�A�R��
�C�?`��1\FM�;�P�as��j���q���Wϱ3V��Q}6w䴒j�����l�l>��xm���	��Q�X�X"ǷK>�c�Y�^o�zY?�<����	Fr8G��|c>�v��#�=p-$��5���]��ރ���t�h�;�])	���C���0��{?���<7���P5�*l����Ǣ�'sK�¼�/�