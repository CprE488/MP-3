XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z�;�u��s��n���҄:������0ɥP�[{}*�ܔ�4��<YTܼ�� �;���qU��yZy�#�ƍ��L$�@�Ј�uE��M���6cS����o�e��? �m����ѐ�o��B:/e�oͲ���5�x����>�i�K"񫋵���� ���&�S�����A
œ���9+8����l���	�	�1q���O��l�k����	���ï��w8��?+ 1�Zi�Y�1p�X~��[�,��� b�~�T�~�a�b%n5�{�v�Dŝ0��=\7�w��y��H#��K��`PI�E���&���F�c��6� sӋ�;"��! -w�2E�7ʒY�aN����O%�>	�����PC�� ��jG6{�p�i{��,�KF|�ȡ ����"��0���}���?�%��w���W��o<#3'?�Mu��y@H�#��b
��u?<5��sAn:�8a��Ч��Nr{&WN� kү�m��K3�̓9��Fd� ?]MA��V��qvנRy�]�L�w��a�Qx+Q�C�m�G獑g�>�d�����3�l�&�P����w/�d��e}�{n~���@.v �[ϼP�� �7�/ЙA���*��]����@9"���th6�D���W/�K��2+�J8=jQ�j�bS\S|���%��-�Y`'�(��0 
� %����fTS�*^2n�֡�s�ɂ��B��'�L�X��5��7��3V�@�4
A���P�C=~.�{XlxVHYEB    2892     bc0��#����k���9У/���������J����o���|������뚩9�����~�쫀OQE8@�����ל��yt����[�V��a jt)xH[�m��V_��������G�%7������A��ZZc�$$�&�2_�C� ��Pb�ǀ�a6�C�*�]��U��j�4�z��tX�.�U��"?5�f ���T�$Mxjo�����t~S[�mAR�cץ�MZ� ���ô�2"B����݆#|l��#���[���S3V]1�	6�mS�A�uT�'E��L�]��Πv"�?�1�����ʻ�翮�h\��1Mz�}�(�@������+�.�������V!�4r�:�7�:*	#U1�˻�>��t� K��[�
�@��o2P��gz��4����qj�8|�鬩��ah�f�^j�?�]\	�.�n\���JE����*^	��о �D�E�Ɯ�T�3�Лo�7\�k�/��q��|6�u�Е�j_�'�o�ʹ����M�w��'��0Ӽ\�:��� ��?4�6���>�r��)|DcG`&C�����S\xzb�)�n��`��ށj�kD�C����/-��5肫�1 �zA��L$�#� (�Ʀ<�b��=M�@���ĈaH�SO�0��f��dĔĶ�ґ�}K̀3l��?W�.t*_��y���s-��$��^��:��k�e�7�#T�nW2��������N�����6#n�v�%t��^�~�7R�4�=)(��Xy�����Br�v
�G�ʴ���P�����5Q�JԾ~�����k��������@�S��'�����ط 4��<R�=�kM�D���8�Z�+�K�&u�֭hf�����+u�񑌡i�7?��(��hl � h?ק�h�^_��Rwr2�ʖ"��)YG��'еQ~�� x����5�b"��y������H�9q��Ѵ��rճI���J���J5fPM[��B;豆Q�:?�w��lJ�_������e�* ���̈́,�\(����b?>d/mm�2¢M�*WGE����t�sȽ�d�w><�Ik|S+{��cD�2e8H�Ȥ,���yyf˜e�b�%!�}ύ�eDQ]v�=�!�<��� kXt���s�Fvĭ�x1x-rRRͼ�U�M�q��<00�>�;���Sb��7���J@���h$�������-��Tp��;��B�o�&��i��1��1L�C�3��£(M�S����U�+����&-Ʒ�R��Q���!`���u�& *�,ѐ�.���$jJW�d4W��6�C�y��B�����amR%&h!�|�ڽ���ӷՁ�n%c�?�J�|Lj�æh9ݶ����d�ڼ)�;X����~̓S���^}����(m�e�uç��?h��s�0�$���6 ��8j��ægh���<m0PJm�o��5�d.�n	`��ns۹���a._�/��ų�E��V{?j�̃[便�s�d8E��w�㍐+�g���z~[�{�7���F��7x�)-v6rt��-䰕�э��%�?��mMZg$�X���4�B�b��iE{M[�k0���3�0e 7w·�z�/�ds59�|�����R'*K�Wɻ��}������D^)�3w�#h?X�8�BI�SaK;�����xKe�R����![Y�H�I�֗�������ЄK���PV�J��i�����n�s�mNλ����ͅ��W��D�n=*i��N]�`8濃g+��?��b8���g[
@�<�ݠ�31<�m��<ls����E�����a�d��ɻ�U�����^���t���>).���d����N7�]��I��}%`�V�3��������I�c`Yzb�.�x������Ǘ)��R��ݫ�I���MY|�N��]A�|KlB�I�c1_�SZps"�X���_c�����/`�U1~_L)���ڇD# L+	?HQX�����,͖���T3G��3�N�����9,��|S��OȫO�c��������m	��:F��lDEW�`
InK�mf1O�U�u!�	t�6��	lُ��&��y�?���ԺD���+��J�u�/T�0��j5/a��ɺ�m�S�<�I���%��<*z���[���p�d!l�H�Dy��8+�[���(�p7����D�ڲ�Ν�u�	���*�=�B@Fa�X����-����.�C� .��D�_�ћV?���Č��1a���]��S���8�ݑ<T��n��|��+�$�&���mH��|��j#I�v];v�c���Ov��������A�<��H�y�%�����18�З�%s�a���Z17�>����y��_�9��z��RQ���r�k�Q�V��ܡ?O}�2�q+��A.�<��k����q�ͅ�!Y�_�M�j�ݾ���b�Q��6��G#6��Y���d���BM�,q�g*3Eў�i��8��m����A5I�9�!��"�3n�px�Qd�S��nf��%Dp'7��6X�<�ȟ�nZ!�C6l���N�D;9��y?	����zN����oE_���t����_٫���y$����~����ܞ�׀D�Q�Ԣ��	�t�]��}�+��[����(L-�NvE/��d4�T�N��М#�|j����9o*y	�<��<�8E��NvZ��?a��q-NR�l5 ��!1��VJ]C%�����
���$\�+ᭌ�KQK��D�q�ET�"��@�.�D
�ۡa��uSh�ij}/�~<-(�H;R��j���-��|���D����9Z��:�o���eY$Tȍ��&#h�/�!	�"��qH��!�E�a�������l_c�\grB�m��<+����2����z �T&y>����ؿ�/9������8�n��v�sȵ���''�d�H���Jb=<��i�v���p�)}