XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��n%�]B��U�6�^���i�}	��*�E�$IK!!~�Ӯ�W&%�q���m�����10�-���GЫ���gp)�,�bEz�^�\%Asd� !/xӭ�����
Y��=���}�n�Wg���@���c<�(�N��W���kB�k/ic�"nI��B)9	�ޙ��އ�!�r�������B�r g�jx��@+FX�5_�Е�U[�$��Я��WL��/9%�:n�"$��ɋo���ю�����@<,>��}�1�dZ�\��Y8��/�7z����Ep3��������8��M?�e��:*�;8׉(�v��3B�:��ycs�GU�kQ(L�"o�#��BYϔ���2�f|k�F�Z���>���[<a��׫ ��{REb�u�3ILXjm��<>����B�]����*�Wt�it:��es�w�"8�%֗4���D��kU�m�%.w�FXOl���#ͫ��C ��n�$�Le���]e)�)�(�:��a;�>1W�Jz��F12�U��@����ҹ�[��<p�E�%#H��sj+5I�$%M��҇ |�$������M��sO@q�Jf~^�1$ǀ ���L�_���9�a��Ha�v��e��vC�9	��D���} ���'];��y�����߫����HU�˕�Ta(���h�'�_��7�n�?۝_!�r��3�j�P�x�nij�uʖV�gH�L��)��1k9!�Z�j���@�������>yx!"ĔPx�\��5*�q(y3Y�(����ʀ\��p}d*s�D-���XlxVHYEB    3a46    1050�-�թF��w��)�:h����v�<`o�d�Cb��lV:;���)ON�YY��#Ff2YOqV\��H���5G��ݓz!�����:5jx=}�% ��N�T��X�s����E�G^>��.����^N�C�k����18��m�����|�1 k3�����>3'��@0�yH��B����������+�0|_*�(�"k��[�. ��	g���9eZui�I���9#]�4�S%~���;d_Y2�ۑ���2�ˮ��ʭ>��lfe�F���8�n���j�'0�D��S�r��P}���/}��X�W�^���5_'p�(�];�*Z��ײ)9MG���~�w���8n���.2j�0�x�-��]���.�J|��\]�����׻-�q��g��ĩZ��=���fR�B��~�4k@P��n�N�e���,H�ef�ۗ΋$�TI�rcn�~���h=�udn��B��R��1�MZ.��h�������2���,��/34&��k�nZI����ׅ����"��4��f���0��h5�;�@��u�C3�Q����:�䡄O�SZ��P����7c�h�J��=�ͫ	Y�MS_Wx2� &W"�l�XZm�_��v�N�[��I�Ya����D�vT����&2D���f����>�T�G�� �:f���6'���G)`wwԉ����;	�T���@%��5C	Ǟ�&i��T�-�7�ǳ�vSS��*Bip�yfv�����W�%>��s�p��͹��B��RZ1r���%��K3p�,[���~�c���I7��=%xr�_�t^\��n0�JJ;���]�'��:��o{7�j5T�)Q;���s�z����ZI����T�&�a��N�,g`:�\YR�i�!e�Rh��������F7�
�DΕ�x�@H�S����cWAȚy�V�1�((����P��3�!kT	?V��@a[J�G"f.O|Pp��X������u��4<(U�l��,�P�̌�i�va]X��V+B*k�M��|.K+��W�#PJ%�4�)���^&�S&�W���"fl�X��Q;��|(7u^��ܪ�C�$�J�)$:3d� 9~({3�I6I�9}Ǥo��D����/++�2d�r�L�oG�Y���2۷�@��B��Ћ�����E���m�4O\A۔�3�5���>P_��������+F��/�ꄢ�dW��y�3{&�c>�@���IE�ǥ0�~�i~��;d6PYm�NC��ֽP�
h=��w���S9%�$M��䊃\�zhYmA����zM:Y��bV�W5�K��vڀ+���P�$�ڷjhM��=j:7ز��F��.J��j��t6��H�X��Ѥ��
���g9�6��7�ɟeg���زR�����8�2~"�X<��zl�I0����-:,��.ܗ)\�D9���ӖXS�L��*EIm�
�u�n�Q���r�4�VR��;Bw�#��kp%N�����5�~��?��-�\dO�N�c׋X�=c�҇��`�S9/�ɾ���0Rp�1w+{��c������N��F1��C+%5�S#j��;e��_ɂ�q��7�c�f�<o2;4k��?�R���3�@(Ac�����5����I�g��kЧ��Ѱ��J�fL]/{ }t$b��X3P����NU��s����mk
d���9��9?���t��䌌�z�3��Pp��t4��jg��J ��DEJ�������^cn���s�g$NR�!��?��K,8�Bz�w��L߮��.M*�i:Y!Sp�C`��@��g;�H5
��qg��s�M}K�rb2^�-���[)�Xh�¾H/�n	���l��F�7pVA��2��Α�@38�1�x�m���!nS���DL���(��	^'pNL� 0\%]�Y��=�-$������؅�%^�b︾�z��k�2�g��@#Ԁ����&_�:����c��J�����T��輀7@�����L��q��ǳLe�˞����E)��J����!�g�����&��7��.mS��S�N�����s���3�Ib�Y�ؓ;[T��X�HH��L��ڹ�{{D&�^���Zh*����|�Tj	��N���i�P�����`۴�
��3�/5<g��x�5mo|9審�m�r��'����r"�7�J�ujnF�&���oΑX��V~�X�*ce�����=ԑ6U�}�s'b"��x��� .����z�e��<��,|��LU] o�ͩx�g�X� =>��5R>,ӆ�뜱~Ŕ�K'IȨ-��8�x.h���ֱ2�&����&�)8�<T}�*t��4�~z�J��T��Y��D�_-ʗTj�$�d�m�i|eB�Dc(��2"܃��Ь8.���8A��{��[{%+���Z��,�K	�� )�uj'P�0Ө�j��F�Kj�U�k�	�V���WQ�u������T�f�Զ8oO+��v��ȴ�KW���s��4G3o�R���赬,�*|.5״���x��ezq���#�(s�tp�K�8�՟�8�6{��^��h��S�ђ��	���k���#NJ�d�7�����T�J~.�ec��{��= D%[�zyC�z$e��~��|w�8�L���ZӬc�����J����*�E�:�������6�H펡�hL��w��59o�����:��f�ᜂ�l��a������(��`N^��>q:���x��j��������H
i��](u��^u����)����*&�[8#� ���gO�ב�
$P{>;�}f �%b=�46��ru��sVNa%2y2⇵|�m��`×/0@kqޘ���'�5���FH�a�B ��TO���� s��5Z��RK4����c�̛,��i:��Tqw�4b(pC��avQv�<���"�ٓ�%��n���z����-`�4h;���W�]T/1�#�9�)T�Ֆg��¯3
3Ij��y����[��?�;�/��E��nYN`(�� �'������2����}�R
��tV>���Q��=�Z���۴Ky� o[�J�r�����mq�����j �y�v�ɷA�@���!&���9�%r^pb�1��~��	�3�}{;�6A�~D�f�ưD��g�:��vڲ�ζ�ͫ�8qȲ��e������"�)N���K��Zh3pO���j�����2�(�˩Zai�;�.�l~�S3k���D�cA�3���0bSWTv�zT�ԫôO�d�9 B�W���d���Ǌ�����:���+���.�T��Q���댶�%R�!po�~��J2O�Z�pJ5$l(2�(��$��c�̐1��bt��FŁ�N�P�I�L�߈\iS��Ƙ�,e<"�v�H�Aۀ?Z�8�:����7���u��q�D�_%���`t�+B	��5��p�\3��:�?�A���j�b��!Ld�]���#d���~�6,���b��tmEs �	��U�v@H�ml%���NFc[RNe��٧�F
~����>j�_Q���q	B��lWʸ�����V��}���41��9D��$?,�"p(���YF����:A�� `��G���͋m?�Uk�Q��&���M�-7ä3a�_���=T?[2y+4�8��u2�{��O<�ųq��?<��;��X��y˯w?�v��N���չ�r���Y�[v��X��	�0������c�Q^��|������H�U4�ƞ �P%��h�a�o���oF�ͫv_X�]ϔ�V�/����~0����_Z�JP��im*��P�;��p��t-�u+���� �z�ߌ��~mda���W��l���$׌娩�!���(�Is��nv�=�?�ڔ�g�M�}�+�����2�1�V�btcb�N2B�����v�k�*��F�2��D�wr���ƕR�HyL�]�AfY؃ �-���n�0ht���uhz� �Y0�b~ȡ/���G��F�蠋SK�D.Э��&Y��O��6���&k�e�Ow�b��#+a���6�nJ<VRYK�4�aLi�]Up�Oj��O䊗�v�?H�����ͳ�#��~���M���I�76�0^��*��dRNy#!;�h��x�>��n�