XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t1�y���>-%�J9��о�f�ƒC��ʈsY4��F�G��@�5~_���N|�`7m��~'�JٵdaN�~��n�3rS@����!�gJ���W�A���
حۜ�s�����@
hǜ�0{P>��6�� AZU8�8�4���S#�&Ů[%��8��lTR�]��ۜ��x_h�B�!�(��f7��TT�\��2�W�b�����̇��`����_kÀ�l��o�Z��6ܙ�P�#�}��g�`-�]�B��|Ԁi��(0U"��5)t����#M�*O���AcJ| Sd3 ��\��H	/#Rzu1r������r/��A�d�%�C�;�(��LE��_=��c󩷲���Y�:�m��Ff�4k��F)�D̀�	s��G��s�|R�-���W�u7Ao8ݕ������V����Dꆈ��
[t�Tz0��l<V#Et�~L�/X0Į��uIu���&oԾ��V#�+؃w��,wzn,ޡR[;ܫ�"����RE��^�7*Ⲓ [M9H^KA��%&�������՜匲ܷ2ɉ�D�UW��x�h.k�R51�3H��"�Ұ.m�.�z���rO}R�%����k��VFn�mV�А�JjIdF ٚ�PQd�����x�f�\����=k�*��歇P��\�{1`0Gh��d�j��;���z�)��c��Ur�m�Fr�M)؃GSP2@W��:3T����@��V{��^"��!h���5v����g5̋�W ��`�Rܗ����
�t���yYw{����n�ϋXlxVHYEB    2892     bc0_��kԡc���I�X�B�,u\�}=T��0��g	��D����������"���Q<Vl6�(�NZR������B}�Etl`�Qѻ~�/v=1=X��)����w�9�=7����l�+���nk�r����9�ˠ�h�F#P��iP��L�C�Ҿ���j��\���w����1o*��5�G����k�o<D���"�޼J���M2es?'1����2߇{6@���蝊��ju�A#-������)$}����Э��� iN�o��z�ʏ�F�'"�u�+'�t�î�pBs��b���=*=�2y�SV�F�d�0����H�KG"�W8����!&�>v8����Af*ߓ��e�vcԄ�\S���%KV�"���s%;%�d� m�!�ϴ"GWaO�g(b�;)Q�U�n+cx�Pog9���U� ���%���Rh��w�.��&Xq����5� + V�0?��Av�Q���N���9���0jn�$����N�.�t�#�K���v�� ˷
�׮���*;�@1w8j>�� Ο�|x�c���n�Se�;-������wM�q�P�Z��������A��]�?��Sf�@�j�u��W� ���3"|��A��PT��&��(�pAb��-o����Ui�?#�r`��F�:��, ����� <�]gdX�u�4�*���Q7r������X"��ܶI#�2=��A�Y(����=�u���l�7FrU]���D��ΚHsݪ��m�\љI��!sT+'�- �\���e�ر��K����T�A��+�ų��>[��ǺH$'��R`/�"NfrD��RT�+ȶ:]j�7����}-y`�����*���
�'��9g�撼�!Z��J��ˣ��!��/��M`=�eI�^����t�J��h8,�8І��a#�e��-)�z�\�
�^����7�;�bR��*�W�+�����$W}oS��j�( 5��si��tx4M�Uwd����a����6Ȧ�C2�+��코ʱ��S��,�͓��-*A�,��)�?݈&���#��:����.e�����eu���P �[��̳���EC{���B��\��2d�{�P-C&�p5�?���A��� ���b�%?>����^��6���}�I�e���b��/�u�A�'�j�+YWV���U�S���3� 󞤂�@nθ�L�]ݯx�	������WԦDTfI�$��� C��+IT��[S�Oo\�ᰪC/�8X��,c["�'�Χ��z3�x��E����{��b�x<��p�б�5���0'�碀�˹�0[�@�Hȯ^ %aS>J����s@OM�&yV3G�NB��~g��U��-���'����lc�)tP=q���d�W|��@�lYS���r	�iψ�Iu���1�w�pé�
ʝ�"UY�Z!�[%�c�J:����f��\�Ź1�ܘK��(�!�.��d�k���r�V�hG�/��΍�c*�VK}�w�`ʝ�~��h��S�dm6�Ƹ��јQ3�q@^���X�Bh�Z0�K�`�Y���d��}W��:G���R���#��nT5C	̀{��/ ��>�G��'�nݖ�����NZ�qc�]�+!������_��p4�� `�+!tJ/
��!�%z�<��B�f�E��`�d�\���3e��5q���$�ѹ·�����* u��//�B߀�`�#I*���` �mf!yn�L!3i�򀣙Ѫ�j<�������SYFb-Ѫ%a�<�De�`��-lOD�؊�*}ӻ]/V�M�9�"�`�S�Jb��s�6)��̎�F��!����[��{b�0�=�&vc"O�ѱT���H�G��zS��X��I�b�p���@�@Jk����'�\,���SX�,���is�,�*�ar��|�.�#x���;�L���<u^=�b?1%h/�x�
Jwȏ��3�)�b< �
	�7:qKlĔG��E��7Z`�˗@h����k8�ME@����a�|�{�C&7>�C�G��%�ˊc/-��E�P�������2����w��0���� �'�QJ��l
��Óy[��ݏ�5Y�5��Ǡk��o�[��\×���Jr��w
,\f���R�%Bf�w�R�8a�K7"�ZtHߨԖ��e�P�7�c���Ls`��8u+���}x�w
H�u}�V����܆��ZN<( @�H���m�5�1�+����5��x-;^Fm��맶���rJ%�j��]o�+66-+תNe[hTV��TVȁpݛD�8�x�?�sGv��,,M|2�)1�L�?E�ZEELe�ٳ_D��V�����ه��&� �D��Ӻ�����a��4�� ���a�&h��(Le��L��HAz-�� ���+@��0�'_a�^���y�q���T�k�!<��?fP��Y��pi�a�DQ!+Ű]�9�g�Y:(��7�u��Q�i�A\�W�u�:"3�+�Z�
_,�`-�G�I�p:�E:�/OuO\�2y���&��N�CO_�]���}ư���<8����c�{�,Ҕ$�n��5���P�S���̓��\����T�Aߒkb<�E.��M�f�D��2<��u᪓}d����l��B��P9s�R�[��b��?5��d y|9��V3S���ׇF��1���2#�ɯ����,k�W��µ�<(ra��嵓�ܪχ;�����0x���B+�c%��d��`M'��1��߳�I�<���9�18Ǜ�D^]����ʋ���-����T�dK5�:�~�ki�����d�B^(#m���6��僓sO^_�|ۄKĕ��c}�<0�J�b�l]�:�'����t�������"Nݿ ��
���o�^��0l�ta+��۷�>Ω%7{Q���}p����|�ݗ��$��=b&F	N��3�`a�|��8�������h�������