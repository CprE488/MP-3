XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/�8y�Fۛ � f�\fH�$�5�7`fQ¯���Z.r�u�Yy�!�����17Y[�h������0U��p�a`*n�f��3w���9�$C���v[����+f"d.""D
���߄z�G�
yJ>�0�W��*�f��4��
�ox�}h����gz�ǅ��8���B�!�@����NXԁMR��{CL��*�|g-�%�?� �rĀ~�[+s,PO;������^��c��k������d�=FF�ݤh޷[i+�R6��������@q�U�4���^�_�.���݀Mb%7	�iZ���/����E�l��)b|t�<��.nR-�]��z�Rh�`��z�?B�X[u���V����ۥO�=���;,}��_ t�*[ۮ��sF���"[;BNŠ�- �؏!�2ۇ�����o~P���76�K䉏u���;��2[_-/����g�{��s�!�دy�s� &�U�|��v��Ko�=I��;ұu���O2d<��Gi>�V�~'��u!�ze3�<�_���t�-���nԮ��1����������q^��"r�4��,��A ��a8B�?0���S�00�V�f�#��&�
*�TA�J���\ĕ��JWY8
���Fx��Ϥ�U��f��ޅ��J�������g<P$�Ĕ� n�o�I���,��v;m�>E$p�����SJӍ�Ip�X^��n�Vx�?�wn������<0:B*���X��/BD����
d.%��r�XlxVHYEB    3b09     f80��mj��Ώ�i�HW�#]�e3{d\��Q}�k���Rmݯ*�j��dI��߾
!ذ\%�og�H�hęQ�dl��JN�%Z�\��o����~�@½h@-je����5�F5дj�-��E-w%����yy�*E��@ҹ�+rP3̻s�"?FΒ����r�#��<�vH`[�+����X�S�e���U�+�8�RRd��&�;?3qR�t�) �$/e[�E�J�?�C�̢��w!�<�Z�g��D�����0:�x���wn\��:�8xO��p�Pf9ol.��/��2ȳ�9��M�Cg"�t�ٶ7AĤ���Ԡ�8��v�aB5�/�5Ӏ؛�����	��bj�v"�t��;��ӧ�L�)��C@�
-��@b��I"b1���j= �!:�W�0���,���ɩw����PG�D�&ڠ��QW�oH/F��j�M����:�ۯ�9������J�j�� 6W�f��� w��+����j)\/�MGf�nƕmE���PLƧ`��Ҡ��_|� ����1���������.�K�L&�/��6+��L	]%$zy�u��u\��R���iy�u+��Ke�,M̮�N�&���bEu��oZ |�H4���Y]"
����I��y�",��
Vo�AzT��g�
�]��jP�@�s���T��&�r��f�5ݑWg�:;����LW!'�u�������w�lʵń���D�)2K�:%��Zn������o�̭�)�W��m�yS�*��I�A�'��-?f�x�-q1A��WBb�7y6�\-?7/��1x�K��ב��U�~���N	����7�jUK��]������DP�����m����r�Y���̪����J�� !UKe?���!�	`� ���q#
7�"�i*�sKπ���U�����,�X�	WU�?~j�.��-���S�8$P���R �����Fr����Q>��cg��䟾7Gzr%WO����_:�?���8�z��a|N�Xj�w��M�����x�N֙����X�|��b��ʴ�����w����B����N �g�JI��'`�����xK�������@����1a�E���M]��c�s/� ۉ��D�^`C���AFA!����	��_�oަEpR��WB�f����_\�P��2����|qAW)�HqV�gwU�@���]`���j�wT&_8˗j����_���x�D�-�`�H��:�2v�XW&����p�Y���[�+΋.*���)yD���0gJ�Kth:�Ue9���zX� $U�����S�9�#���߰ܧ�%�gp��Ƴ㝭_���܂���a���k"��R�p�Ee�s.�{2u�Il�|�5�uE����a\��5�1�>y3�/�O6S_�X ��\*����|(�� ��X�߬6�A+�8qc�l7�����+��)��[G�J�!Ѝ��j�<���Yb?XTt_L-��*8������`ۥh��i7Cq�������G�n$��H3V�Xy�6����/��W��
��ٍ* ��v�V�t��������� ���г}�.B��A�����b\"y�jR
[�B:��g�+��!R�����3{m��!Н��َA������ͣe��ԳuE�~�6-寺��]?z�����9��a�9�gL���k�ƻ�[��e@�%�;�^��BH'��� 6N�8�}��	! $�&�O��`�֡��X��ɡ����]���c�\c�u'}Ҙ{�lK1Ǿ.��E�K8�t+�}-�� ;���iu�ⅸ��|�&�'�oƉ����*���y��y�D�|穋$���/����i�ܝY�+�.om'؇��e�?�ؤ*�2K(��h�{���@�6a�j��G�z��9��� ���vn�<���L�K�}$�m���6d�p2����֔`�k��'Pް�&G:$[�à����ʦ�BJL:�F�S�J�;��Ǵ��� �X���2!Dȶ�'�d}�G�W�+#�<�5"�� �e`\�z���]����]d�se�V�t�F���a�]�T��5�?�b#���b�-Z�z?F��:��D�5*��
o$>iǦ��4����l��v���(�B �YGY�3�&է��0�J&�jT�f��M����c������u�B�	̸բ'm�fb�*�U�̾�$@�5Pv����_���xF�W�s�����U͐qS�=�䣮NA�6`*h�⚼�d*��������`)Q�P�D�b�;�%$?�A	2~��f���^�TY�������l�~^�5�#e@����/JQ���j	Ʀ���)g*��,D�̰I��B�\�.�ҿ��~�R�N���@�M�`b���l�ɭeY�P����-���m����[��F����}�����v>�����7��rW�'T�6��M��8����e�2��%p_�C	9�9�%�G��Ɲ��9������
�!p�p�45�	�0�I�o��/�(�_wr,*�q\�KQ�N���O3V�QOv;'�GS_��E�oW�o|~���i,3����y)�E ��"����!�!�Bp�����jc��4b@���CpJ@�
�1&Y�]�T^Cw�
"j/�m�d�?���G�N�������9���1&�9g:����K��R�sSb��J��3�ي@z�&Y�X�0�Q���t:G�ث˘(��8�0|E���&N���G�4냼�8����2�S+y����aB�%O\(�<(\��2�"��kG3�e/�R�8~��>�je{�ŏt�@eZ/�T|�m��m%$	/'��� �ʵׯ������e��!�q�1m���@Gg��.x���W�,zT�}�V����@����o�R
*U��M��G�zU7��#ɛ��f*�_���Wc\7�x��s�'՛�;kȢ��a�2��iyն�O���V��9�a�y9��d]/Z�(���fо�c�ˍ�4|!�o��:�R�
xh<�����W;z@��,B�ǖf���!�$~g:�@^�`_�����{�	qȲ���r�����e7S9�i�r�?5��~Ť%��]!w'��y���P� p5D��u�j�����)Ex�ݩ�0�eM:7���JDJ�<�3�C+��E&q������ v?{1��1��FK���M/f�ǁ7+�-���C�D���#�6�~�����{�
+��M�$�g�p��&D��
�yҹ�#n����v�A^{�L����5��14�<=wK�hBTԢ�|pF?���{(m.rིᙻ�/���s�5�cga�����)&��.�ت�o�f���'�@�'�jaAmR����A���B>��^#m;�K�qzE�vܫ|Bч���9.��jE�%z�s����@S�h��K}���������ܛ�ёzvp;*��s۶�B�ሪ�,�	�Ŝ��G�0�������<:��B�c	~��'w�*�L?)���@v����s�%�l�]�:��V�(@j.�I���yo)F������7t8Z�ؖ�a`bb7/i_��`�=Az��N6I����:Ձ���^E�>J�44���MSg<���ӳ^��8a�����z�Z�I8.^����̫��:'.�r���\�e֍���Pk在1����"�ǔ0У�W��,N���O�@e@��oq^�8#�68�S���v��q"2"���˿��18NFqJDl�2�3�%E��&j�ӗ�������ω����ҝ�w
��E�B"1:�\���\�	8��m��4$�7�_[o��l�O��8��x��6D���Ʊ7������M�������%�~�F/�yM��ܹ�]�`�����4ojq.���2+Fs%t|���.'4��Z��M�7���Wj�Oy���X�>�Cbׁ�