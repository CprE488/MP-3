XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���s�h��4V��L'���#>�&�@�n~�Nӹ؇�[S"t,{�Ug�S�T�&�V�U_�[Slae��#-�C�u���#i[n�;����+E*�}�1�'�r ��<[�9�����>\]�4s���H��b�$@iNk�.�^]���I�%���v�[e���P�r�I�-�����o���%{ċ��N��As��H��]�S�Ӥ9ZwA���svI^�y`J�ҋ҄�uD�=��+��X�㠋Z2LGWF? ���m��a�5�=a�(�>�s���.���N�"�X\�Z��}Q6se_�ʼsX��b3�$�I�@Hj��ֲURH�L߲<���r%�)��~�g�@��b�h���J�.�؁4�a��?vC��o�|T��7�����,�u?3BV��j�9��+4�5ӎ�|�X�\��([�'�������$Ƅ��20�m���=<�"�湖?�n�3�{V���^�oi�\XRûֻ��@ᷠQ5���M��mt��Hc`�'&&��)'S��fjHNӄ��&�L�(91���)o�Y�Q�r^�ŐGق�`��h����XE� 6,�
;�@��	Th��r������(j_��6`
Lr�X���s�}WL}U���;`_i�Qe3N�` tC���>]ط��+��YR(�/n�ƣ�9=T�.n��[� ��[��6���J��"|6�I��%�"����o*���|�z��ؙ������Q=�p�4T�?�a�x"5����6�9XlxVHYEB    1847     900�q�O?��!uz���-Hl	܉�΁��Jy��n�u$��9g��ycc�q����䰼�يԖ��w�.*G?Ĝ0����/����*#a�{فFON�q��r|��*����� �S���<-U�|�*����5o�ۆy��#�S�m�~,�E�B4��y�� ���-��f�D�#1K�\�KF
�Fc��8���Z&JI�D�-5l~mi����MԦ)��Rf��=,}+����x�����_n=�81���j�1��!c�Z�y&�������L�}��05o0�| �|&&\-�� �y��3���I�.�]˒����~����_!8����r\����)��;����0&4����0Q����r5\~���̘�'����GK-K,������\^%�x֙��iY<��ߌsfQZ�NbU�w;�� �h��@E�Q $�C��_V��;���G��,a:Bmw�8Y��:}Z�TA�ɯ�-�����ɳ�Û	:����Qo"�<��2����V��Q�&<Ƣw�E��&�GJ��B hW�(	&He@
R�Y[��.��$�(-�c,b�N~E��/�F�C٣����CSP������b�&���}'��S�I��S�R]�|���@h9���6'b�����������Ԏ��(iY�
�M		��{a0���-V~洀qp�!�
���%�"�r���`%��ɂ��t�To�t���w{�z=d�����T��g.4!=����aqt:�e ��"���*�z�I�f�!K"0-�����5)K��4lޭ��;���XM��A]R|K�R���x:τ�UKӸB���Q�!u~f����9�����Pi���Vf��QK:��o�x�1��Ib���u��l�W���e�N��;A�5�EēN��|!P�Cf��o'M�qڱ&��~���
��2M}ɲ�&S޺�N��2.
�l���>O��ZO�����4�gÙlU<��[�b��t�F��!�(Dz)��K����lONN$=�r��D�aa�O��A�T��ɑ ���ZV4��ͯ�5�td,��?#�.�D�n��7�u�|��U��<���`!Cv:G'/�cE�Pöi�qh~:���Q�����h��)�V�h�uq�G8�)\��G�U1����.�q �����������kD��p�[�< tR�i�l|S�9'���L�vD��<_N�G�'��>*�Q�E�w+f[�\;�!�/Py��~BoMLջ%Z*0 �7��tgd�F�����9cFd�:c��z��Q���$�U��T�.7Ѹ��EB����Ba�ʙЖd?c]KLuBbB1�&:\f��Z���a���yҩ����%��c���Ct�xR]ѽ�ԥ
I��&�ϟ���Νf��=�ru�-X]"����\�Z�ȗ� ~f�<ufNh�b=�%�1�cq����?݅�C�Ẍ́X���h-���s�]w��P�J>�����Ҷ4�:# �"(���
ŐGݎ�j�v|3���NZX�b��nx��<��jo�{�/�%�.�Xf�E
�G�k�sY���qd�V��]�2��r*<���K�����a�n�p��}�%N���	��*� �*t�!R��n��
$G�z���nD��}��u��\�*�����Q���$ٸ��WGuGк�m̫�����:Ȃ2<����{߲�UZ�X���6GQ����,��<�H��ggOێ��j�����ҠI�3�/eWJ��{����"�3��P�n�/��p�YA�� \�D�7�������Wm��-�R�D�ڤ�d5�I�x�˜q#�%��*�^j��b��@�Ѥ �Nl�3�O]-pi�'6�Z�O��@�vP*�`�g]����ˤ1�"W��`E��l��=�o��Ҧ�tk���~.=l���''�'�Í��U�/2v�p�&.�����e�Ն�I�635^B̊�VM�z�p����Ejg?EJ�A�M�o��#~ֹ=R]���DP[M�����\��V:E3TQ�Zt�,��~��}�&7�Љ�j�
�cղ�mb�7���m�2B����sr��f��L��n�?��z�s�}JG0(���Ĝp�/ݫ0����+1ј=��)1S�!y�͕(#�/��q\�{�����!��gL"���~@@�,��/�2���Z_qk͞'<�8W(�*8m�A]ʭ蕀��u�,�ʱ2�Ϲ?���ό�GT�w}���4s9L����e6d�,	-PN���ͯ��c-Vi�P��r�P۞Z���α
��8��H_~��|
A���X