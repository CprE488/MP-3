XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����;�D��B�Am�[7�r�	��&@±�9��]�EyF�A`�s˒2�lĸU�*�d���ε΢ܒ�!����o�N0 ����P'9���q_8�Bvո�/5f��6�s���[�ҝZ��vM'"P�g����sV���ϰ�#���i;V�w�����$gA��V�.��!i�,	2�<��4�>şz^�#5bLP�Kc�W9�4�5,���������p4�볩�-�r	s�����.]8uPz�R��B���I�������{��}I�Kl~�=SF��Ț��>3���N�KQ�v�U`��V>�~ ���B�6	�9�d5���J��]�B}�֌�*�TI���X����]��"��s�;�-E��J��,���,�zoj��2-�B���}��\x\N�1���M�`�e�������x��O����b�^*��vo��w�u�2�RYg٨pTBn����s�Y�dk���o�@��c�݀,�`���= H�!s�h�J��<-w�G�<����@v{��<�����p9*D˔z^��K�B��v�=AD��u��W�|�& �˕2s�����l�%1E�;��t>��3C�W$p�,C�X�|�R�,��'|�haʀ�u�tJ��a_�>����xO� ב�N�%������?�c-��q=�f,�-p��� Ē<4�cw�I͋zlKqԢ�|����@�)Is`@���:���&� ��ޯ���^��ZOS��[��w�p�k2Q��.!�j�N���P�B�G<8����gýB�X�\۹XlxVHYEB    5224    1740�ͦ�r���g~�L>]s�r�,���
y���oyķ�N^5f�hV�o=[�(�ZO�yOO����]Z!�5��T:��� �Z@&v�M޸I����ʎ{b����|�W^ܥ-P�6�l����������섡��'Յ"hr�L�V�ĭE.�%�J��O{T�hj[��K����F��6�=��A;ȼ�T�������7��^�}��Hs��b`~3٥����IU�~����N�G����m�>mb���~���[9�,7$�ڲ�c�E+V,ϵ�tS�[���/�r�s�,2��!J�BD��� 
���	p\ЫQ���6��c��L�	�4#�7���trQn���wF��46��{J�b�#E�|1�!K���k���=}q.��DQR��I�|��F��X����/�-9f|�4L�����col#����V�sѶ�q'�y�����#���
�G��w��J����A=�2Z�,�k)���e���M��+{��sy��Dӥs�K;�=�YB��~l�5kk��]�_ub����$�rA!J�-��_��G�G|Ƒ 
Ќ��hrK�>�o��s=�I� '�N�;J���Q�A��32�l�^${�2�C�BK:�G����[n�rwNo�V�ޕ�&�|J�閸����d�Q��fLx6��*@�����;N(�6���t���<�
�)g�k�+�K��<H�-�',�����/�
��nUI!r]��ӯ�����<z�?� �1t��ܒV*���!�ȬѷǇO'�9�R��
�}]��M�\�k\�C������_M�K�~��O8�w��u�2��2�i��H�2�r�޻hdr�U^_6�z_�W��߇���(��C��(��П��X:{�\��1	 v��$�M�p�ydԻ���������7/`<(W*Ue(��I���^uCM��A:��Ɠ�`oAs[�X�+��Q�9>����,;��և�E���(BS���a>��Y ٻ��UZG�E 8"5��QQwe�^�Q�[������W>��ڌ �&���!DP�WH��&�zt�D� @LG�<���<�> �}�w鿡;��*~��URtЖE*2y�Q����"�H�S��p�q��V4�I�+�Sǚ'��2��Z]9��}���x��N���bz�G�q4����`-G��;�K���	���u����c7{ʴg���IXq�����]�Q3�p
�w9�fwkb9�*�5ɨ�6Dq�m�2!�<@�N4��y��w=��V�e�7�me�:�`��y�������[�7@�� ��q�->�/Q�P���_�Wb >�EN�]�^A�nR���h1�Q�	dA�L.�>��=���$/��/StAV|�h&������y��y��#(���хBso�5U�H"��/��}��RH�i���M� �G~�9C0�=�Bs��T�7퍺q<EG��ǲ�Bh��=�˼%>^���£�����i�h�CT��+�R�ٺ���d�@b!�ekl%���V���XrSv��x���	�M����^J�a/����+����E���
�����S7lқ���Q��E;�z�� d#�D�_D��@�;�[��:�����S^��-��<�X-C�pt�Q�c��?lԛ�P%�Æ`��3���:��ֆ��Kj�y�A6���=�K����c6M��"���lY&�e�j���pu"8�f�<�n	�6DPh��d|�n��_|�c2���Eq} "x�b�p�x9R7CxxH�6��D�SW�L�/�7�����H��V�S�����1�>��3:�g�iZڤQ��N������`�C��J�����=�N�R�gV�W�f���4�5�,�[��$���> ���ɳ�o�^c��5��5�	�_�;����4I�T���8zQὃe˗�����Ʈ��~�����=�1Ʊ9̈���;��&��� FŚt��ON�d��zM�D�q�&bh��8u�2x��"&IQ��]�H�7,�zF�1_}38�몟�bXw��ʲ��9WN��� ?fP���^Y[�OLT6;��3Dި�t��u��}��F��utr���C����>�	�t�nAp�#���a��VWl�L�:H�&���`ؒ����3������e�0���$�U؏"��7��i<��.�97�w���PDF�R|�it<xϑpq4{̨��(�|d݇�#N��.���ZNjk�-η�zT�����tMĒlr�>	�v�&�ߐB���(h��� x��jn��xMV�������wycc62R��K׶J+A�`-��ֻm���-�oX2sQܴ8[*��>/P�2��;e<�����@w^a',����E�꫞l��i�'������k>�L\NÚ�pl!.W�"3������/�fq³��ip����T�V ���lr,����A
��!�����jR=\��<�j
��z-�[����%�]iX9u;>Fm���h��Hn��^�m9 ��S�&\v���жL9!(�
g�Ow���o2c���_�1��k�Ow^�2P�\
G�9VV�W�u�z��к���
���/�(��8tv��$hm�S(��&�'Y�;8���)���c|MŤ�� �U��/���Τ����J|2BB`�1j/�6=*�A߶O�P5�߱��lq�v�o{b�H��Ӵ���Hw�kK�:	9���R�ob��uU�t(��c4t��T�A�O0�����`�X&
A-5�Ql�B!�̠� �7�u?�)䩸�ǚ�w��W�ko�c��v�G`s����ļ ��� �8�y]Q�/MG=�,�M݂�yn"*��%��x�>|�)�o@�5,W��<�o]؄���N5p��Q��/��mA0^ҿ�)s�>M>����� �	-> "���(̹`��Ǫr��,��x?����ge	���#�7V�G]�R��U�����i{^���ַ�
M��~.��z�w '�֠�sS��5껟1�z���D��`�;H�߷�����_g�39G�y��/��~�ϊ���@�D1��H�OB�1c��P{�x=�*���O���5����%�H:�~�m���AK�-�n�
켥㷥�rŜ���X��W�j�e߭�tp��&p���������E��^d�Vn4��Bw2:��{���6'�7�����˖��/���(1gz[x��ܪ�ʞ��#��m`#����]o�PaC�|��E"壿�J�e����s�:�/������6�a������ Y��KB���^�c�dd�ֳ{P�EdQkk_�)��A7ĎNBU-�����w�Ꞿ�fY�_I�@�SiW6��ܧ�jQI�+������\s�%5E�X1S�(��6H�q���7�$��cܬ�J��`{�Ǧm���w��?,�j�����󰭳�/Y�	M��vF�^�M��D�ɱF$��P�g�������g��rذt'�Dl���7��T�a�Gw�ؖ�U���;���d�u�κ�~���7��.{-����va�㡢�������qe��p߯$	{�x���WI?*+-�i��@b�����DOxS�F�� �e�#�+�6Ĺ�i����"B!��mg-�]��.�yqm��s)
	�I�$��Q�`�.����U����%���fq;�%^d��z#|�~�_�A�p��k���X�1��,W�K�~��0RP�(��z��l�/�D��� �.L�����v�_�*ǁe���"��O�}u� h�XAR�w�(����-�����T��L�}�_Zx֨�_\�&?ì�AjPGw�9�lT�"��Vr��l��
q|[ջ�����iXf�I��"�Q�����z��_�̎u��nk"\2Rq3�]=>v�;4��{H�L2؂��̆z�Nc�x��6}��� `��a�3���2�����xl��$L�5,�Ji�k ����I����a����ӎ�W�rA� �78,���e3������go��f�&�(E3�-�ײ$O@f�8�)��_�۸�H	�,�[�Y�d�;����}�:���lz G熫`�jx�&�#c7���9�&����4�c
L7��9g"�._�k�ݗ�Lx����C�wf#��ž87x����#)�����y�x��N�
�/|����(�T�R2��������� s+ߖU��ӯhn���0&��B�s��z�}��X�Z���ynS�4��8zЈ7�i��Qu��F���WO����5�M���/M�,�I����G�Cy�Q��2)����D�H`\�N��x�Yyi�@�R/�y ܱLnʢr2�Vķ#@��sz�B#�X�)��0�z>!<�v=�������Ԣ�h��l��6wI��u��C��=+}���x�-�VB~���]��s���{�OV�)�&�wQ�\�Ѳ��.f�9�j�%bok������}�QIx^�U��5~�dH)T���#:�.���)�{��,T�Ѐb��.]�A_�PDs�p��f��Y�[�&+�- �@B4�~��Ĝ� $z���d��D�n�&��y}N�ã�U9����1��s���`4���Un�1~H���/wK��<k<1|㖰�}�H�5�-HR�̔��	wIn�<W1pM�آ�;�C(��p5����ս�"d,
yč�k� ��
E��2*���dj���46�+k���B��+x�C�R��'��y��'z��Y"� p�82�����1fd�	�1���#1�Q�G�����hU&%�7z�I:���u�?�<8��![L�+r��K��-�SK�JI0�#�ϡ����9���j���M��l@�Ud���2��Q1u�`��#��
�^Ldj!IX��T�:����A]ث/{�i�t>
��v��w@5-%TH�JE�Ѫ��X�;IO�8.�>�=���_�.\��y2'`��ڑ6���J���Qc&+��a8����M/��>M�����)�;�MQ^����:)��IG�F�ׅ!t�jG��XT���e
%E�C���J�� 2�''B�MC�35��w����$T
j(�a���Cտo#iǋ�<Տ��ꒊ������,�9mQxF��a{�`�S{�8~�/� G�^��?���ntغ��
dk6QWWFQ���S�Ů�{���b��2ӈ"��N8���k�爘m১�? ��+�R�NX~f�dCyK�$����t��wR`�;B�ؔ�+\?"\��KO�>L���X��b�T���f�}�7�����rPB��9�����",�a]E���O�`K�m�E~�=h����E�~c�/��y�����4�p����39%�'[�$�<�V��/"Bl�� �������8~��ѱ�4lD���!��B8�g�Q�d��SCu �Y�h%�����?|Q_�i�S�`Zs��k��38���bi|�Ρl���H��h*b�4Y�|���p@^��:��/z���kcߓE��7��7 l����ƊŸ����i��>s�a|��6dK����t]��A[�.�����D�Xۺ�6�Ǝ�f���b��!�����;��^y���ڟ����[�Z蟁{'���A!.��7j�o�R�vP�m�k�e}�w�i�E%��#�z��ג��~2��w�{$#Uer��.��c:���W��,���3�DB���#+�,��x�����i<<��Zvx�.NӴ�g 0��֊���m�^�ܤM�u:Y�@�,o���q��u��<���Y^���؀�9�i&�� .}�O�h0�Nb����T��[L�gl"����
̙��B���d�r�E	bG&�7�N��m`W