XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������?VBFZ��qK-A���*����h����BUEӴ���X��R|v$� !�D����X�Zh�>����������w�%ٖ0��k�O\�%���VD9�)�5�-�@�f�v���8�-�D��]��z���R��he�S	CP��.�L������1)w�*�E����"��[�UU�R	0�i�-�`���{a�4B��*��tU�Gϵ���bO��b1������;䒆(��y���`Q�K�F����3�t�/�b��;�&��T7�989��xm�P�iD�ʏ�-��Z��//��+U5��WD��e�M��Ďtׯ� ���A�'�c�X�f�v=oH���v|dKӁq��h=;�ףs�k��@-��t��=cr��R8F�_��M�Z��R�u2�����˒��M�o	��cSb�|�ɩL���t�жw&!����˾��z�>P�
$+�_GYcY�����w2��9f��^	&�4��!&Vx�P�c_e�v�L|fE<c-`�:2�z@~�<����5n�5�;��JAZw=a�^���^c�Q�����1j=�r���O�f��brż��0�~fg�y�D��G�����&�����g�~b��W\%�j�wr�ASH�����yO8Pp�qo��S�^-�ŝ�,9� � 4�c
�?P�
�ޤ	��b�Ϊ��m9`���L?b�%��=������hH	��wUZ�(���!O%�7	fI���r!zڿ���XlxVHYEB    2b75     cd0C�GYw�0�!xS�$#��̅�U�}A�6�!^W�8�2t@��/= `�N]�I�r+B�+���T�x�E:?I��rŹN:0o���پ71`����=�暛=j}*oN?�$@E�y�5�v�6�:cY�DM�Q��*4e���;Q>��۲��M�#D�f��e��!�rN�:"�����4@����  �f��t�nz/��پ�a�}�(	��	��j��0e��Y��T�ZJ�O�unǜ�?���.� ��5/�̋Z������z�����  ,�r*ފqգ_;�$�9�]�=����s���k�����b��O��D�hD�����Ȏ|�S��(?�&��#<�.�����0���sd��"���W�C�09F��7#�O�0~kz���n�������09ѭv�`�d��B:���2U%��{�D�~��Ez�;Д�w�qJ^�.�[S���vi>G$��5Ҝ�'��l�2qJ����;�_ײ��p�y�l�g������sV('+���R|�]8��5?n�)��8u`~y�dU9�kP}�W�n�R�q�1��4B4_������7{k*�1ѿ=0���j�H;!]��? RM$������0A�3�kGھܜ<3J��ˌ@����[���T�I�.4-d���o00�I��nm�JF�io^ �����rZ9���� &X��p��������k0B��c��ח�5ns�ͱ��,!��N�M�Աwu3n8��w�n�_��X�z�s5��\����h2U�0� �����ͯPn�׏H$�p��R����]e���5 �Rz��9/vf\G�M=ڧfԣ�l�]����q�/�0B��������
G�p��9���T�|���.���!��R����L��6ԃ�#���|����J��f�'.���GU�m�2����ҩ��6䩈L�=��_��TT�Q]�y�+K8�wh�����L��8R���,��K	�*�#;M���`?���o,حCW*
2bg�����q��Wqf�5}��  :r��}�ݎ���r�/�w���""D�9��Kp�R�}:Ǘ#<�g��>��� ,��*N��<��]Dp�3o�5������/���s_�(�<��%�p釥챔d���lr0|P�FvM{.gM����*�VA�[�7��%�%ht����ok�!����726��2UVѱ5��t�j
_�{�<�c#����Hj����%>�ȯ�f����2:wji.�B7��>666�%��f��(�	1�:��u���t��t�t�����Z r�ˋu��y�`V8s�񓸄�F�u�|5��tRfQ�&s2Q�-��7�#c�$e���<Z%v����y��p�1*"�!P���@��ޘ�;xM�s��.v�
�ݝ~&� �M��t3�H?E�{	P��=�6LX�4E����SV�P���w��J��CW�g�x�L�*8o��2� �|�)��gv���:��j�� lV�(���e8��
��������?�u���W�#�.��أ��#�$���cHП�D��w����#�d�hY9X�|)����$r��RU6�$�+׮�n�@��I�nĪ�׺�o�7�tBN_����c2�r3Uפ�V��Y���4��{0C��K�}�8�Q�֢j@ubn����(��r��Z�cS�%��YP��%�����S��;(���d��Wp����J�H�\��(��(�"�p>�n�@,Q�)�)e�@}�բ �]e����1�@�ynwʅ���_#����}�E���W=i�$�7*�\'���a,���Y�#�l�e寕�+����eG��џdTo~ 1��Vw{U��A��b������(��흢I��:�V���m;8�l�V���a�\��?�y��������k���S����p9�+w���O�]8_�Y�>&�Fs�.�����{z��T��q�����o��]�sׄ�"�L]�º�?S�ݡ���w��Ɠ�����a	��h4��%�}�Nt��\v[2q3Ǧÿ~��Aj8z���.�ط:n��p����$��s�`�+=S�`�
=lj�c>�9ۊO8�}�j�*PZ� ��2m�U����o�y�8`%���vV���$Y�FPY��`�|xU�?!d����<
�?0��Fcs7bz����4�B��V��:�֒/$�X��y:;�+Y�V��1���a�Զ>�H�4�m�E����7�-r���q�����9�[� �C�b,����~؟�ߨe�[��Rt�Sx�g_}M΃���+3R/�(�K0U:�&��h	"Ĕ��{΍[��B��6u�r��I�fC������J5˩��t��(��aR-!�X����'����Ký�\+*<�� ���W�K��yZFż�av2���o��h@�����+G�f$P �7��#ܚ0>>���	�� ג���Q���#��=O�JH `����� ��o�1���r���^�ڠn'��t�%G|o��K �A����¶6�g���7ܽw1���w����}ׁ\�2���/X^�+>X�GmG$	��l�S��eY�)v�s�K [nqgZ-�n��.=��# ���HF$1�����6Ӿ�O{H�H��-Ѫ݁"�%�O��H�o��uЕ��N%�X����i0�@�I���J����f�0i@���q���!B�$�!~dى�I�	l�zi����q�E^����1k�^��A�i��?9â>������lb[ݍ{����4�M4�CiJ�X�� ^�	��Vpx�s�,�0aٛ�h[py�u�h��02����!ޅ�PZ��k�?5ӱ���N� ���~�&�F�SYl{1-ܴl�C�ggY^�bSp�Cs<��m��a�Ѧ��e< C�;��������_�kU���Aa�z����?n���AI]i�_��b���������멶���g���>�_���0��>4q�h�/;���4���<�\�'Y�!	/��smݯ�X��F4==� ���y���dS�X��l��)$_�x�Ze��������ׯ�4��RT�|�ߎ$L����;땂�ݽ2'�!�p�����N��'Ay���T8��S�p������c��C�3�@W���c
�E��s�g<s!���Eȥ�x�O������{mi����EC����}ψG�iS��5C��)NZ���B]�K��m��`�����y�}���j>y���Čӄo��Ϯt,��a�X	�m@�(��H��VJ�	