XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��N�}���>�l�0׹�v���F���d�/c�0>����{c T6��*W�fL���nw&p~�����v���kgGV�i�����n�:.�����7<g4���#��ȧ�	�-ŏ'��rI>>�4�Z���f���9����
�31��C7��9�kOL��{�%���vXo�}�-���ڲ7}��{R�n�(�B�pY�,�:.��*+��>���D�I˟\�<�4���+#��1�%�7)L:�eу��e�+g�L�<��]6��Cm�O3U#9�#�ĊL��-��2����,�}ҎoC`�K�dه��U�0}�a��NR�κq�օ��)�_y���_��~����	����{���N�P��>LA)i�	O]�>o�T܀ M1�~��h���7�ۯ�1*3/0V�3��|`xd���P�<
�Y�O3�Q�G��A�"�6͡[_6�Q�W���'�]۪I	?��Z�O;;�*W�������%�Ya���p7�I<�/�,��iT��E��=*�V���8�ר�ٟi2�qR8
���s90+䕃(0D���/N�5B����>�`��_���r�=�O�zE$�Ί���
I��S}�i���F&cn��~��X�u懓1�mN�x{��0q�:�
����0w�`@�� S�q]>��"�;x�d~/��~��MP9���*�����
DVE�u�rz�R����/`�+*k3Ñ���m���Hl��)1ҽ��J��m;b�;w�m�H���hFXlxVHYEB    1ea4     920 �x���X�^Kg��|b��.�
��
h_K�J$��h�:R�r�+��\g�[:1Gf�=�X��Vf\%�	� �Z���-(� 5��E椼�����pJ����E��E���k2�Q�X�PTW�z%E��]]�F���R'� ��I��w6	�4�>f���7o^��i2L�Z��6p:�j���O#���oUT��?0w~����y]U�Ǘ��(��������V��'����:�)}��RUrĆ�Ҵ+��n�^ٍ��\�9���m��8�p�����/���j� J�/��8n�}N�i%i3�X|w���tL����:�S��:q.(�����ۣ� �D�4�YE,e��}HU/�NM�q�Ӝ�5��@nN�빻T�&��}{0p���!۠O��x��>Q������������G��-��:� lr��Z�w(D�c�6�!5�'���i����+��޶(��W��.׭��-�}���X{���.	!��:�C�|ŝ��K��nZ·���N�1wU���h�#=ނ���į�#b��t�VWQ�|~���<�aNo,n��.��U߸��<*�G�\UZd����[��02 Ñ;�b�������r�[p0\�I3|;�B/Y�zz�,%��
��vj��{9̶cƎ� ͲC����B8�i��Wv��"��q�D�/LRc�o��[O���P�C��V�f-�p/��,��"���Z�P��E~,״uQ(�m���P|�J�q#A�G[8�y'+��k�ٯeT
�?hD5�9C�$|�MՌ�	0��:�o�<�> �ՙV�U`�����Q�i�"��$��B{������e�����.��@�w���+��b�s����t��aa�A��������Ж�nx��ʀ��f���	��B��B����;����t������>6�qC|�*�,"��*���d��X��!ig��w�"pB�.������6c���G���T��f�%mT�J�k:ɰMlJU�AeGW�X#�*���.3i�?���X��f8tZ�CV��:I{뺵��Y~
N�yL�z��o��0�q�T֏U�|Mf��/��A�}P�F:Ț!�_t��I�h��ʗoz �!�g��ƕ�I(�k`��4���q;~���d�^�E�h�k�Z���Yܚ1')Z�*�9�~�� YF��Ӧ2Eo;%���~�pL^^�О��Pqxܵ����u�r�Q�lc�+��Q7{ ���H���c8��ԣp�y�u`�Aú��7��9/��-�Af�Ϸc�P�K*I)�h_$��􀆁& ���pD,�`�|I4)��w,���H$pP�Q_��9x[q��O�g���r�W�8�n̽���庢1#�X�G�l����3��{+�6b�@D���Wg��d4?�:�8�Uϣ���'�$K��>���$��X�^wkA���_Ni*QbO���"$ލ?�����qO?׵����
G3�O��x@C�~�]	���6�;3X�3k�^�`<�9Vp�>ظ�7�+M7������Z	�^B�u��K�_���i��#�I���S^�%u�ț?՛99
D�vG�]�Zۿ����I��N�do������k�o��_Y�����o�GvOwHs7��C�m�������K�v���W=�k�򙏄�zt꿯�`>?lR��':> ���
��>{I^�~"j=�T/P!�;'��<���+�w�6BHi��<k�Y�x��QԐ.`�����P]�llO~�����ԧ2�l�󧚄�`wj�𱂧��[\�ܣ��`�vBrg��KPF��wۧ)��tR4W�n��<ꕓ�O�i�Y��U�J��т��oM�_P�瘍���)QOX<\�)&�d�0���픤��`m� �·��H����y�0�*�[=�2������W�w6emHgD�{�wI�ۄ�R��CoCr!�@��ֺ
�=5��[��I��r@8x�=�-&R��O5Ö��m|ܒ�d�f:�mm��Vf#Q\c�/���T��GU�+j`���[s���~��&b��,|n'iYz��W�钖ݹ�K,�]	%,���x6�9�T}	�U�z����q�$%�S��`�X�́��K������ j5��)��i����qI��_�n�Xƀd�[4�P��Mw>X�,9�i��lթC��L�x�O�2���3�N�:G��|�>25���ABX}칈$y��Ip�<���廓!2ſ֑���;��7��8��tyv�~Q"���E�?uy�q��s��d��u!�a�4
V�|�Jˋ<�ő��8ܲ�����8��v~)����9����