XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������ƶ����z�4?�o���Ii��A?-:���Q�P���z[�|1���A����Ek W�|�|��1=Z���A�:b�0���_'R�n��>5u����m���G\�'=�H[�M]Xd��sO�ێ���}����U��B���eKpb��9R[l��O�V"I15*����z�`��a�p��u
)b�#�t>�Xߧ�B9pj�<Q�j9H���d����0R9l����u�7C}�>+C54���q���� 
����qs���+h�A��o43��I���u}���,@� m�_v�PgM>�Rd�q6��bux@�{@�sd)���@8�s����7Zfd�8������t)�P��2�	�;�,��l��Ծ��u�����bp�Xi���U�|X��6��{ ���]�B�s���g���4�����fe��5�T7��H�YѨ!^r,��qǐ&�Q�.�AM�w֤sE~ 蚓�V���DC��Y�� ЇB�W��dI}0k<킊�����hpct�KQ^�$��C���Ҹs�\�vF��ȫ<�!�(Vc���C�ʆ�H�A?�aSƈ�h���:�u4�8:8凹7���9a�C�Vn+5�ctw���<��^��}�ٍ^���������Tm9��F�G�z*����k;���
���xl	4�s�@���b�'��-�C�����&WZ������ �z8�:s}h�@�H�OW\e�C O�q1~L��~c`xׅdXlxVHYEB    3da6     fb0��v�����r=��a�s��^�g��6v�T;l�bK�D3U�;���~�o��Bs���a�z��A����l�g�Kθ1�`9,1�������XO"��6���XLf`Mlr
eR�6���	o���Ԅ3�&�>�[%�o�xbbt�����i0Z�a���|SJ�X1s�_iE)��RN=��\�?Y7���-LfC���Ua�Sv�p̀ݐu߯��_�'##�C��#i�o��7�Y&��>��I�,b�Sh���Ç��FT7����WҌ� �����ve?{4\z>�#��v\&9d�+��
A�7k樬�����d�^�,[P��t)h��&7�7/;lr[���c`{UA0I�=9�e��ec'�,������~0��U�:�֗�D�G��|Ɓ�u>ˣֱe�Oؐ}�+��
$кEL�n|��o�\��"#%�Όn����s�q�(��!��\���a���D���}��Z�S��?�.e��\u��&6Z �W�{VzӒ��	U���4��=�����&0����uءT��n!u*��{�TH)��� 'K.K.�6(#��x�xJ�s�@e'D�,��O�W��
�WӐb� 2�"0dO� ���>��;��B���G4��	���8S�ߍb��=�IT�@��;I+-�,zT�MW��Q3�J+X�쿑�l�!�o���W]G��c܅���U�~5\x�͢����;�&�Zi��8Vv.�㵙�c_�.^m�m�ض
y�5"g�|�?��&��]��5nⳙ+,����6�5˧��垒�K<6��A�:���;��E e��zXډ̽��d`O ���Ƿo�=��Tm��0��^ˡ �j�rHz�7�-���ީt-㱬�ݼ�3�2�Đv?X�7�dr��:Ǡ׊ȋc]?�YHi�zU{ � ���Ɍ�t2Gƈ��3!H��� �"�,\��p��.�D].^�/cfeF��@�`U���۵5�_��-w�Ir�-J�~�ZE핽�?�+��`�U!�L�"qvg��>E��4�U�E@�?)�&U�N���G%!7�ʡ~4TǄ�������Y5f�&�s~�H��1�Z�3Pz(�Q�3Ӡ߷i_�B����$�Gzc��������sXU_��LM��K-qh�O;�S&�@_��J&���(ƅ-�'N�d�Q��,�N �ݛ��'�X�@ʞ/P�Zi�v�ܼ�xD�Z�f�=�	�F䴿j:*�RJ��Y;�z%o��ڵ,DR�

q�>�D0��,��z���-�v:�՛��4����#�t��e{���`���hZ�}�G��"̚���0���P�W�P� ��9��O�R*(1��,gԀ˳��r?Y�AwF��^\�w�#��bd�,�~O�p��ș� �rp����[�������₺�#>$QPtM	6.m�)ɧH/h��KD;�jc�'J��4E�w��xq�vʱ��d��<�?�ܳ�_�7ݣ=d�/©��B��5�"�3Q�WTM�5�H�S���J�#ZQ�o
6(Mcآ��U�ǫ���4#g�V�y`�F���%ɽI�����8(����p,�ſ�R�.����q�y�j������a�,Y$㚞�0��S�9�$4�D^�yb�u�RGm!*OŬv��!���{0L�J����P��B�(�)p*٣gH:����a{��v�f�<�b=Fx���9gV�"��s�G/R-��U�%!Õ`h���_*��)< h�N�^+
�ADM�얊����N%	�,6���z�`���;6�`UYk���]3{8���%� S'E�<��~"E�v���/\�hoГn���'��s�=)g@H�:���N�&�>Ih��L��� �U]J��/͗�!�-_�kAt� )���<�B��d\�S��Y�V���K�_�s�̓{F�`5
��TΑ�q|�	y!y?=|P�8����;��8U0�we�
���ltZŒ���3R���l��q�OU��sr�%Ã	�`��%����mX���V+���&D�Q�^@�� Ȗz>V�������E;�d��.�y����Aq�|^����d@��2e���H��p�u�K���c2�0I\L
/�Jqw9ct���ʦ�0�Z.s���v�S���{���p�$��·����RV�\Z�?�2�Yb��	&�w9�&b�?�J/Lq@	��KK<|��MUv�[Z�O�"�Q��iiXUL{��Fc��xhA��t�����xWv��4�d]�(&�I$���Y�Lt�;��</��"ʮ���4�2u�{�BC����"}yQY��&u�miH�"�G�'Z�M�3S�)=�W���=�?N��@\�s��X��-qtY�v��t!��8q��͌4�mT`\�f#�ƌ�B.2\��(�PC�/���ԶY���N��n0��Q�'�&ػ�?����lo��lN2�S$�*�OR?�Ij��e���n�T����;�U'a�����t+p���Þi�����[v�Лo|;Ϻy�H��ע�9�3X�iZ�K��?E�J~6)x����K�&,���Lߩt�i?cٗ�s-a��/]�@�m[B�1��"�Y^+�^\.%#�5AZ� ;ǧ��d����_��ih7Ub��gE�nT��ަDA�v�Π�#SX�)���#���ؚ�5��@8��ȅ�s�}P��|�~�³�s=����T�w�E�ۢ�R�i�EFwi��C`h����	�"����U�pF<���'����b��-8�d�P4����;�4'p��1��ݜ�Y�@���5�p����h{��4��C#�N��1�T�@Ȳ~Y^_K�����r���xI@O�� �M�J�PNd��>�\L�g�����N���[�
����m%�1`�_���g�?��
N�����I>�����ƕ�T"�oǱ�b
r�MOE;8	q��녏j�irG�Y�v��^�CA�3�H% q�n���K�Ե���[�+��f���b�
�sJ��ԏZ������-�5�?�:���\	 u�g��\�}2L����e��WV9HH��M�ϟm��֋xb���1)_O��x�g�3��u��K�hiǹ��߷��v��*Ϋr�A�qL1���"�Q�B���=ZZ����!�xA�@�0�l�	�Z����H���T��}��ғ�v��? �������]���a��_u?&F���;���"�u�&�2	�6�5{����'���r�����=�˼���o�j��U-�]�i�7�˲�C\�����mWɞ�̵b�˄ւ�c��WA��г-�KĤ�R��~n=�9Ŋ4��_�_�c)]������[⍋�P��<3j���-���+)SZ�k�;��h��U!_���*SW��w٦)��d��ȷ�dc�̣8X��0��?I`bL@�s��T��^=�����+���οf�LtI���"�/10s��se�G�?�0�S(CA,��@w���V�e�V΃��"W�7󝚀[��}���:Mf�w�`��+Aw0��&_�ڰ#9�I/;��y%�$	W��t��z��c�U���-�
/�/�K�T���k���q����)�5a!�bB�d|8>�(�� \"�-��Ƕ-����=���KEE9I{�㝭W������\���/�\���"��Y�
^^\���嬜F�޿���)1.�5�����ƷI���*��V�������p���.Q�R�T�HO�j+1{@uh��p�
�e4��9��DT��fcu2�����6�1�N�S:qQ+.�<m��5DX^e���7�6����2A�ʉ�k�V� '�m�E��
��s!�!,���U32�j����'��3���ϹL��o>��������K�?�V��:�t!��ϱ��16D�6s��a�L�Zӧ�~���꽌ǂ�M޻�6�S��g��4��9�+�6��\��~�X�K���̀��x��x7�: