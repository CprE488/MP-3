XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����5|9$;�����ѳ*��r���U�Xad�ow��֏�����#��.�פ=ɟ8�#��޻�Y��*`R$Nk��e�-ͺ��FM�0�[���w������.o��C�0��ߩ��y0w��Rօ�hq�X�v��kɌgw���܀�V�/�U*X-�K8�o~,��ȥ<p ~���m2CF�i;K�7���)~���R^&WֹБ���7$u�T�TW��+�Yc�s�����!	x����I)����£�e�c�Z���S��b�xAX[.����W�޹�<���M"O�VV ���"��@��FѮj�P�Y��	M`�"��u�zX!I9!�:$�����s���ϲ�)�U�NHO���-!��jϒS��l:,��3��u�c����Zj��&��cI�
��>�SL5C�$0*�:q�2c��RO�پ�Хz(�%�6�4�A�ٔ'�)���n�y�������@�JU[�gxK	k}bFGNK.���l��>���'��\YuEK���/��2"�.檭Icgw�@�i g��$� ������>MI)-���A�-����5�K����Z�]}���0>Ea؎�3��3y��bB�����۹��Z?\���d4�L��H6���[{�#y�S�s�l#��o��B�۟[D�����;>I�1*����ނ�C
@X�K���j��s�}[�����F�{D��,{���z�(K:;F-�g݁�TçêM[�k��wH��!�=Z\a�M P��]۳XlxVHYEB    5866    1100��)�9�=�ߤ�����g���^�W�ZG�`����<�������kԦ?��6J!��rd&d����!���]E�Od���
!�ߪnj�ͱ��oGA��Q����?d`(��C-�UɌ,2���V? ��1��ᨅZB^�(�\2c~>�-Tß&�ې4R ��3ߐtzt<}�+%�U4¹�wmy,�5�.��"�$������߯��[��j�W�`�����5sM�-lWs��t�@K��$�4���������'3/�����=[�YI�@�8����N��IN��e��CЋ���du0��7ܯ�=`�1W��|�A6�D�!�w/�F�~ޯ�BU�C`i=x��.C���`��5Vi��ie�a�;�[�Gp���u촓i i޺�S`O�rL�#Eg�{R��]��f�W���t�U�yS�hk�x6�������Qz3�TԒn�0%�<��	��pK]�j���Hn �2',�N��&;!���;�d��Q���
�5��`Yc$�r^�����%ub�'�Y���7�+į�~.�,�Y�SN)�{ʶrN�¯�}��M$�F��FQ�`�+��!��aA:.�jtJE�l��&�i<%B1X�nŪ�Oi�"VKR����=7�/AP"��XV����l�1I%V����A�0�)ܱ�A�yj}W��J���k6"��T^w��^V ��Q��V9��K�'���E�l2uc���U��!�)�1;o6_����f�;�+���m�q+��,�u2 ���ڀtd�<tQ�B��@�^8�?R|vg�E�7�K(�e����/����i$�B�C��pt���m��z}�z}oy���=�L�.�Pcl�
^�(�`��su�=2|vK4�m�	lT�JD]���*һe`�7�T�(c|��U��]y6&�]��@<	A�6�i
�_,(6��_�\ɴ�X+�Q�EAHu�Ls��A�L��������^�A}@ڳ�"c�/��Z���W����A��P(JRX����fkM�a��q�κ
AVD����+O��|��Ko��c��q.?y�BiÖ�^z��2�d�W�,M�s�����4�:��\�/��gܾ��	�G��B5iTLt��l$�!�v��o> ��1*&��ǽ�r>ߠC�J�%9�L7~�i8��ki���E���Z��qt�I���}�ZF�h̓P��bDxN�ɾG֐s�f�7��L�E�����>�5Y��u�.���G�}�������]eF�{�I�Q���]��m��o=���qme���g �XZ&1�['.M�]�������j�00��e��t�����?�HܯKc��9�GD���p���?<A�]�0��&J
���c�^�2�I =p#�Kh���)�(,�Ca��K5�&FC_2o�t7�cd�@9���4D70�ngW���h����g�<���vv<S\�
#�@`t��Ův+?0����{&9��p��g �G^p�$�m25�e���{����e:|ʕ�r��u��<G��冻ni�g���N���	�ԒQ��$ >'�C�V;Y�Ku�&�ZXv�$J$N��� �+��-�{�9d����>��/K�~O�m���Ӿ�U���8���y��s�/c��L�Ĝ�u���买�%E�y�w�Ʋ�Ef��j�c4p�X�čMz����[ ܼ?s��AsU������q�S֧�{p�9�� \ޫ��y����q�K�� ����2���B����ڬ���'�� ��L��v�Lr��A�Q��P�E\,������ʳ��K� x������9�@�;��%������'.�;�j�՝|�[�m�%������F��"���J��`�,u��$��t+X�2k�M�;^>���E�ԙPI�߻�v���Nj�٤dpl��/�k-���}�w	]o������e��dl!Bџ���V�0��<�Xg���B��<~�Όp��;?�ٱ�.u7��d�<���2M3��|�j��>_�>�h\�ff�\�Ik�[�z��)4�]rW�Fl48�����K>��F���H��ʯXAi�	���[6���Q������b���6�Y�u֮�姣:jg��sH ���o��gM��Y���|��j���]���	�p�4�s˱�]�a�����QU�/���l}�a�kj�Qd�T�h�d�m���6�I�(� (��q1]W�Y�DMm�����ϧ��$кlN����"�� ���r��x��L�>�xT��e�t2�ڌ��������!� ����Ǖ��ˇ� ���{­���i�y��	��8����X�f�;�TE�c��c�6���+3_p���}5Ք�e:U���4��x#r �{S�@h���{4���K#:܃z�j�W��c8�?Gb�M5� ��~[�fYZ��3E�x��rT���!��0��tX��z=ui�(j4�)(��A���Z������Ny��5a��y���]�̿49{�oB����$V@�[���j�w�V8�og�Ƈn��Ut\�޹pW�@�'H_+L���˱��`kjV��es_�ďx0`l*F�\�� <�l�m��I�!0�y�&�Zg�����}g�d�гMf�5D�Dgꗖ�m��K�ϻ������[?�?4;3UQ0���R��O�ٖ�*5�	Cթ�]x;�ndr��*yH�����~b"�_�r[@C��=ӯM�B����#�x±/��	�hh��o�v�!H�E�XĐZ�8�_�b�㯌
z;'�Eٻ�Bj^`?��k��Wժ�@?2=�d�,���A�9D.>9Y�ior�<��Xg7�־F����w.͜O~KE�S�<EK���rI����+7P�B����ى��-4���<���Mc~���>X�z���[1�N'ő��30�J/Y�d6A1���+�yr�Q��JlU��j)�W�گ�Y˓�E�nĄ��+��z ���m��ٻiZ�5�H����-"�e-%����wǌa~z����ҟ��w���zz*�e�,�i�&U������V�B��fɖ���ǆ���HjX8o������<-e�h� ���C�g�pXr�㛃J�
�1@��ͨ���v�f�ŞE�°��)`�s�����28��[Y� 4���x`7�C=N�w�����٬����L��9:����__�6cų�VL��m\���-O����y� ��|�����0��}��D�3Nx����ߗ�D�5�MR)��Ix_�YWq������KT�1=0t��'������E��ȼ�%�p�t6jṑhH��^��+���d9+���j !z
΃Le��ma
�z��6�ִ�#��%|775͋g�v��!sT�"Td���,×�CN�(#�	ن�/�6�s��k�6��W]6Znka��ZAnF`�O�Dmҭn�����ц�MQ�<VJPG\g��� A���JG�xVA���x�1^����Y��e��0e]��?�`P��2D�����j�F�n����I�4Թq�t�
)sG��Z����
��~�.�Os��xw��Wٞ/uvD@�,����V�uD�L���m+v8gJT��M �����r�B��#ph7�����y8��/7_	�"gbO�=�JO���G�'�Ȣ�QR^�)��W������4��cP�M��7c ��S
"��J+�u'i��M�L-Vs
�LBf�їm����\�sM�
��ZW�eT�@V�0?�hE�9H��k�4��ENX[�G�'�4�l�ʬ� 8@��"a����K��]�Ů��Q����/8�`r@��?�s�tY�ǔ ;�=����W`���bWʗ(B��oL-X��������w�h���p���o�mA2��C5e\E�)o��&�������Y��e"��:t�#�+�14S9������
��ԥ)}<B��#_� J\�7L"�F
+d���_2����e��ǩ$_�3������qkԜ�����<n�R�����G�٬�5�n���-�2��� �_���jMoe2��x�`I�!����jY���Ͳ�9p��":SK�릛efh�C56�k�8ȃ��>�aH�&���� �-T���{�f�"��p���|#��֖r�������C�v,y�+�}��;,}�k��<)]��U����]�G��_��,�+ozc�+�����	L�GRv6��H��ڵSK��NcICv�s��HKȶ�P������!L��dzl��J,�L�(%��Ν܉2���2ˍC�6U;�Ѕ�R_*bw�