XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��s4�! ��@��6�x!`�i�?��mB��|��I�������t}&���)�7YZ��3��3U�_v����U#mr�{a2z�}G�~<Fnπ�X���t/r���L>�ĺ�sZ4��@���c\i<Q�.J��{n"�#�8���JζyY:�0�%#�;P%�����3c��P�LPi�a��7�d~c�PЮ}~�ĝ���\R��%4y#|Y7s����%x�p��S���������)����=�"���$m�8�l��L[\�+KNB��y���}�{��T�i��gH�>x����z�<{��@G�4K�{�:*�?�3�#4�����:H4�a�T�/����ac��;�>�;���:�{���HS��R��8���j���PQS\��ۿ�?=L�$��w_�A�Kk\�I�RϨ�&=c56n��B�1�E[��ÿ'<2�[źD�	5�)���{�a�E�	�ŏ?����$ܩ���'s���u��]Y����'ܷ鸖��|�l۶���Fo;�K�>��+��X�'lyÉ�r�5�zH� �'TЎT=)*��M��}y�R"�}~� Vw�%S�Ь縇43eE��V|փ]���k-�t�׺�[?���T��W!po�`��d�t���d�O+K �9<��k��+�������������b}֝6E����f�d�w9�*�Βs��gkr�n�<�S�0�>����(E@7���4��U����f���9����L�����n4g�f_L��XlxVHYEB    2326     980�Ҧd��=+������O�����a��]��,��~
��>(d��S��&�0~Xo�^�z��dⱬI�I���
����\��)-�>?5��*Qk֓���m�	^�'-��� m�Q�����������G;@��5��1�mDbu�I����U�:�����k�Q!x4�[�����R�(� 9�/�z�6�׭���N��Jx� *�?8���&+W�_;B�@��8n�S	�BE�ljx{F�\uyPj>������
� �5��|
�㏏`����8f�|���l|"Ϯ�'mw�}ߵVl�V"N��C��r��rd�;
�Ɖu�*	���t �k1�<|?}&Bi����6��ZA�"N"��3�V3�J�Uj�8�2�f~���_(����I4�G����u��@�Zc�=�U�b�����	HJ��ǓmP��W��Á�=	N�C@W�4�Y�ǅҸE�C/^/�b0�<�Q�K��8w��F�$��.�	T�L�_� 2<����u�1�&%,�Tq��b
��}�l���#8�@٭m��oZ��)K#IR�c1wN$W�G(=�d��G����*R�+��r�O[�
�^�^��UԪ�� 5�N�p��1�̯ Q��#g���@�JǤ����>� �w�}��fV���h�M8M[�����򜈲��o;XC�c4�6�H�t���'��l���o	A�@"k�O��*B�C�8V2����z��FJ�荷��^�̈́� �Q����Q�J�{<A�t��m�cF5D!��%�_ř�}��!f�=N�:p���m�MZ��W��|w�c���I�+'��u�UJÎ� L����X8�9~�O ?կ�#$�Fu�'�֊�\M{�:3�B4��u��z�m&�g�A�R�ш�*L(�na�ǗG��Z���U�[T����%��s����ӫ���̧�����B1�}���Q�5,�ʤ�X�����L�U�R#E,+����Ƴˣv�1pHt�m�)r�3��A�8�z�`�wj��ےW��c_sB�>����rv6b�%'F ���"rf���&	��i����c�z��^��9@��ioEc ]rm���I�l�rw�Y��������v�=�6[9n��3�����|���r>T�Yc����t���2�v;�h�K�V��£�?M������2�����2�tՈ�k�h�:R~f��$��'Tg�Y�x2�Y�M��������������ܐ�pS�7<Ѹ�l?w^r	�����;�AR����Tr�zk�P5��(qb�U�^Pp��*J���=N��x|�g���+?��ޡ½b����Ě-X�	F_6 ���F�)�g��RS�����mXG�D��%~I��������Xফ� ��Q-m� s�9�G�}��$?�F��y�ݕ�q�&/�J��/8��m�+��4ؗ_�F��j����pC�?���FR�L�
�>n�z�׻RJ�����N_�!�S͋����.C%�ׂ�N���R>{1�}�2��:.�cIlU?]�Q���� ��=���th<ܹڭS�Ⴁ8���ə�\m�R���T���)���϶�;?L���xW��^ER�L�c6�W��:>�r7ǳ�N��L�_^����`�s�b:��+B�R+����:��w>aK�m�{V��K�^��W�X�l �WLv��'�֊=�
1#���\�m�����A���b�He�����:H��t��{x�m0��?�Q��Ur�{r���;��@�h?ɒ�#�-�  I��s�L�u>ُ8��(�f���J~	��MOW1GWL����i��'�{�0D��+>��� �u�L�V�d�lt�^��@��t�x͔q�h��)��@�I{���;�x��v�sw�y|V�cm�g��L5��k��Q��"��T�<M�B���/9����q$���k��� �'m����;B+:�ݷ�Ir/�;"��zR� ״GglZ�1���*�0�D��Hk�`�}�.cVY���<U��^l�n��7�a_"���M��;��%M7� M D��1!�I|(��G��溬
BJw{�Ѻ��>_���Ħt�sE����,���y�]�͕U���ʛ_D�2B��g��#'��G[�ΓO8F�'<W<S�!������x����Ҽ1�ʌ�ܲ�t��]	S/%�߅�P�1�X�:j&��B��E!h�_�7r�0���ZOѶ�b��poU?��(��=ҁ^q2P�ZF�B��J?�dN��p������2]]��=�K�G��
�e�{�v�(ƮSvG��|��D,��&?����[T����:M=�Σ���8�$m<����{q�٘�la��B!]���D6�o�+���h�M?&��ܮ^�4,7�h9R�J-��W�� ��Y��a~����̞@mJ��w��"