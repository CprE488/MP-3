XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��e���^���^3�Z�(���3�L��x-���j�����C�%Z�_,4GzM�*.#h���_C=�tF�ƭK�*^�����\!�D�mnޣH��U���#��@�ᐣ�|p�فE���0�IU�u�УV���胀��o�n��<�'���B�UY=Nkr��8�%K�oA�H�c�˻��|VQ�{���)��.Y����L1�(���^�E����_h�+�������-RM/��/;&~:ϲ�p�Lަ�v梁�����M����*`V�/c�D�Gh^	ٛ_yI	h�����Nf"MS5��sj�U�EB��f<lF�m&���8�ǁ���G�;�#+�T�4}@T�A��0q�[9"�%���lԧOY�K#�)H������S��C�N��O��~+T�*
P��x�`*t*l�$@�:��p9�&3�:���'Fr"�~c �R��x+lb`�#6���ɏ�]�>_���vjZ�Q��6��e+I��.u������"~kӟ���g������	��kу�W�s9�?��uU��:[�G<[n�NGO[BB�g�p��C�~(�Z)&���V~#5k�������|��Fo"iV�ژdvnN��$�� 3.=�[��$\��z��ey������<g?1�im�!L���ژd�+sP��K!��Ҁ+��v� ��	�x�+nƷ��7�W:�PG�'����;�z�ϫ�-�\mBӧp�rk�]���@�(�S�%/A���琳J��M�N|��jXlxVHYEB     e07     680����9�rY�s].�)'�����B"H�d�,=�l�����p�����]�:���s��p;�%7KB�S��2�[�=�?G�&pR36&;.G�XZ%{q'e�6�+���i�E�yʬʔq��/ �J��'�����ca�V�w�EА>�&�u;E���`�����aD��yu������M�[RZWi3�@_S�9pE{w���6w_LD(c���ѧ�	�%�7���U΍׺5)U(Q@v��ܓ.�ya��WR���=��v���
���U��q��+HI���_L�����m﬜�벺guG;s��rf�)fu<Z��BS���E!I{zd"��I}�</s����ʝ^�N�V(�r���f���e��+
s�n��9D�P�8���������	���7>�>髧9ڎ�5�2����1�w���6��9Rg��[�e��-���b�`�ڵ0���e���#��f�"�Rk��:�0��/I��Yr��}��Rc�%b+t
K�������^`齏��*�	է䠧 ���2"W�f7�
-�5��Y��e�t,���T�]1�,��XM�pj�tR�����4�_ s�î���K4xQ�%����F�^T��������/������v<6�D�-�/�r�6�_'�r:!q����8�LNd11?:�O�#wU=�Xm�>��ȹgO��t���#��[]bX����75"*l�F<a>	��Ủ�[��o�B��\����qn9�mZ�y�cc������W�I�$��6�ϡ�U��2��#1͞?����G��[9=�J#�B=�kk�~�{��#�2M�����vخqI���j�A._�Gmן�s�L�sd���LE��Qe�#�W�h����H���9#4��w��N�	�x������
5�g�����&R�D�w��fUh�ސ ���u=H�]f�\\�%�|�x(��Gp:a���|�/��k�xӝ�`=5����{͠h`�
���h���5w)>���&�1��JB ��U���	Q�;���� Ohi;$��-����7�$�u��/e��f%)���$�4a��c���q`>8y�Z��Y��Z�'�[{�$�߉��-37�c�˵�À�'\�'�	\4�����@�-3J��*F�QF�k��	)}��)񜙁P���5?�G�y��x����MWwРK-������b��VJ$���B���H�X4n:?�K��A ��Hh�����5�����▥�[�p]Q`�
S��KIt12����1��ʐ����B��3�V�P�l[�+/6�&ѵ��N����gt�8_)�&BG�S;Z��[l7P�;�����L�$��b�7Q��z����M���-�RP��5�~����Q�'E)"����a���'EU�Y1�L�����＃�`dxs�d��������"��s��G}$-e������>�p��M�l7�:H{m�E���:2+�B#��!u'X�:�_�u�����K����$Q36�1����L=�~`�r�w������'��UϷ�}bK��OD�{�
ܬ:oikRK����x��F��HWS�)��&����uIR��'PR@��ge�MNFM���8��o|���e�Hhm�,�Bşp�