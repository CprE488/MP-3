XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w�xѴ��MX�ģ+B���R�L:#8v�zzغR��:�{[	ϤMR���\�����
�3�X��y¥K��6���w1='���s�H1�ll���a0�V���v'��@��o�j�Vkr�(KX�cl:U��0�0�b�#��6���S�CB�]k�sU���z�Ę ��W�+-�H(� 0��L�֓	�3�#v��Mj<�
�!l$�{��`[ڃ�s�01pE!'7���j�)�9�^�;oj����k�bx%<�dP��Pg�b�	��#H��=sZG��3�M�y����������f�)͠ҮG��=U�x̲�=g���%�o��=��eY��F���������lP��>� �l�۬��1��e�zR-PK;`�{^,Bff�t ��!�w^;L�m�Uv��D/�C�}��<�3� r�"wv�?�W�$D�\G����-ї.r��=�B��i�Q�Sw��ش�4~en:��_�Wo���$����ZA9� ��,�U�J����x�Y�hz�M�ȑ�d���Ob�̬%�����R�?~�����-w#�5�c?���˞)�Sag�B*��L�����i�MQEߺ���?�;QО�V����VN�q��N��,F�^L�����yuf������=
�!�����%����-��S��?���R�Y2�9�Ջ��JG�cM�{�fÙ_ºF���IVw�)Y�R�35��i��͊Y��nw�^�H�n�j �XlxVHYEB    da59    2e30jxY��x
�ؐ��T� ���,Y��w;�X�ٺ���O Xē�TZg~�f�d	�o��]���E�l�#E��Nϭ�!��3��ZQ�m�b-�.E����B��`w�WƉW~|h�=�]X��E�t�3w�����!�nFO�����b��u�r3R�ư�.}���=�5�YH�x�� �.z��ul����U�\��������d���'����Ey��{=�q$.��*�]��ĤG(�v��"v�6���m)z��gMr2�㿵H�K_,j~��DBl���x�-�qz�n�ו8���o}܌��g8MZ{�W�^���2׀$qq���=3O �K����uH��S�{ ��v���D�h�dM�b�*�` �
So�:����q� ��t�=���$�yT�ɏ�ߨ�q��>φq���ښ�{9�*p�P$S3Jf��9f�(Oi4)�3�4���2�v;�9BJ[h�#��Z*s?�����D��y�{@:@�/��0���동}��\�PoW�ݐ,ߣ_"�ҧp��e=E��$7���Y��W`�W����%i��J�˻��u��S�^L����t�Ϗ���D�������g� �2�w��v�{�м7��$ԛX��E�D�ջR���_�����b��C��	hL:A�[�M-$�5j*^��"g���W̚�I��·�s'�5��u�^��bm���L�%�E��l��5�������_��ky7����r؄�������p�bwMh�����W���hXS\Nؠ�L���7F����k�<�ބ�qv酫��d�=��f	�mh�Ɨ;py�Dn���<��n��+X$jߚ\��;6�X��a��m�*�o���:Z���묷@�c���Bk�dxb�>�v��&J���蘿m�ׄU/�/����N�������";%�eS��%�3�x���2��٢�t�y��"J!AeM�?�ȣcЛS�&Ϳ1����@7q�j|^�.�X�Q� ε���P�k�@��˄k9HQ���`S~��3k;���@$S��(4�d��3��g��<�� ��h��%!�#�%�w_l��uZR�t�c[��T���ۮ�����՟�P� R{2� ��8i��R�c	�м��G�棆�E��U�a��)T�f�ڝ�W%+0�y?�]�Mz�-ъ�����8���wnXʓii�o���������Y k�Ymr����f��_�}I���8�m\�w�R͂(�7�yӼb����3�����d�f~��IR ���4cV[(�rI���G��S9\d��~]�Ԟ������-���
:�G��m�����X=�K��P�8���j.@�WW7���\$C�^�Y�p�oǵ�a�/p_-���֠���^UgM��F2��햵^^�mH����.e����64P�1^T�k)��G�&��'<X�I���=[|��p�4��� �nx�����? k�`>�u_��ó���飨���3�$9���\5�7�7�j
��Kux�z1��ҵ�Ϝ�$�1^�E'���	�|��pIZ9ͤ�x`��[{��X-�'�*;�cjB0�j��߿X .�B��Ţ��p}���ƭ�Z��O��I��k%��׎�F���L�슱�?���y!�4�I4�=�4��I�v�k��
���g7��u���۱�}.������I���ݠ�(��ATo�c&���������pf"�E��L�G��||�`�]c��N�}���B�6��D[1���R4
�tH1cɕ�$��>�@�ƆR�U�Xx����n�c��9�2��ֽ�Fm���G�0'�FU��RTkͨ� 4qM�߳�N
��'��1<���u�1��jU%C�5���r�}���Mj�5��j��t2Z?��=���3]@�~�)X���w�x��@M�\�+��kP��2n`(���Vzk/��A(�Z,0�C�<czz<��) l�d��RZ����s=q�����-DJ�ƿ(d�Fi��]u(#ȋ�+�/�zΒ��k��ܡ3S�,s�Mo���!%]��Â�xM�$�7����ɞB�*��|;�� 8t������ʩ�_: d��c �HQ�1��!i��Ѩ�ĝDc���g|�k�K=ϿIKZ>������6����oo�'�RF�(&�ҳ��ӕA���a �j�k��V>7V���ÌVd����ߢ�0(�D�^������*��9Ċ�-*@H����L��}��d��= �_���ٞ���c�@�V�$fks#����b귳��Q�m0�.�R�L. -���2�he���an����d�`n$��y�����a*L+pXP�m>[n�a��R$��_[��cO���҄�`��C~�e�e RQE�h�l�mY�@� N���C6mX�l�C��ެ8�Z�gv��F~��?m��;X���O��E�gwɊ� D�C��r���z� #oiE���6ߑ�^Go���br*`Nܷ"�����2l�̻�"e���j�"95���]�i��Ǩ,�	�'��y E�K��� :���lۦ�=t��q�E�����q��*XEJ��e�gZ�:�M;y�"9�Jy����k�n����^*h�+R���[�#�}���S�`#�e#�/(ѫ���f\#54�ͳù�n_�$O��رN8��%4yx�a�$�~ׅ?��h�,yL�(��ǥȹ}�'l�E�|�S�����u��9�w4�>�ϰ����Dh���������i�t�(�J�r�x2h�����&x�/\_+�xw�;�(�Ϥ3��"]	b������\*��o�� :V�����FA'��N�🕨�k�xt��C��������o�R�J�À�R�B
|Iz²p)4s�@*��@tM\�	��>�J���������P�1��xq�籫����sy�t������x�
{ͫ��ko�hB� ����n�}��X�����\g۱�ݻ	�����C]�s�ׂ� ;!�&����:�j�m�	��e��)��v��&�VQ�����T=P��n�:"�8̈́t}�Hǯ��C*�)�� �� ��{n�������3���Ly�z��[�ސ� �bڟ�m�vb�2r[����*���Nx@�<�Ru�	k�DYb�`�F!��鰕*��EFT��)-�?g*�	y��z;�CӒ�]!XiyJ���r^a��O�?��c����:��=��_L�]� ;����K�FW2V��94�\C]�᜹�إ=���/Г������wv�(�*+
�b��A��Q���"�o��bΆ�Z��|`[LY�HX�!:piВ��
ۑ'���Rm�m��[�#F�GU����<���W�5�	xL:�BMT:	:]�.�U3ܭ^0%M�L)W"��T4�����|�п�ܬz�|�!o5��Q'����])"���E[瑶����X�����4�>ŶRwov��I/a�^�B�>VT��(»�4��_��"X�`�\Ig�B#�'dh)����=�`u��d~vY���܁��'�n�qc9Ja��� �*���|�@᎞�Y<����A}��+ۅ��."�i�J&g�bƣvhk���d/���+x,��."D������u�1n`a��7z���G����������4�w$����]OZ!Ì�O�Qeɱܱ#S
����i�!b��<Wn;������S��xн}v��t&b!�����+�	�A��ݻw��O	�c=���\jfMƲ*iIa#�Oz�e�5�|%2)J�9�#����z���|�}��ej�Q�S˫�,������K�/���i���MƄ��ԉ���@�K��G�պ D��L�-��I����r�@��͑�!���u�שE���4㋮a������l���a�=�w���͕@�J*/�K�Od:���S����]'b���Av�Tl�9-���KT�.;��~�F b_�J��<�d���ϻ�xa"��Ffl n�|~ޣ�^�X�����*�k-�l�FA�l��9�xe�{C<4w�J��}WXɏ�����C����Y�� �:$x�y�(���C�ܪ�h�mM	��x�T^d0��&,�F��5�����$�^�W,�!l�����nߞ�䃮�ܱ�&(l�0��K�Z�� ���A��-��[S�n�M#�I(�;�S�V̸��g�|���W4���N��m�Sx�}G��9�/mI���xʎ���vs*�E�遃�B�wX�36�C��#���E[�*���a�[�*�������y6%��&B�%ĉSz3(9V�ݲ*ԏ$Н��%���� �K�o6#���f���;�Vn^��x{�H��y*�E�s'3���)Ƙ�4.D�[<��{�7�~����=7�x�+��˔��R5�?���r�=jۂe�9ڽy���p��s+�c6��f����d[	q�`����h��z��y?\ؔ-t.Id�
���
��-�j�m�ou�ڱd��h辞�lL-�;��ʦ�i\�ZT?��
TM���z�ںYHbF���!#��&�-�K=�PùY@j6����Zr�ႵXɜ�$���;A���6?yO{��8v$����glW��WO��ȣm� '�ê|oj��Y��v��	lU��%˺|�0'g %� xN3%luJ(�Yu{�y�a,R鑛���gM~��(8�=}�z�cr���osә�゙],�n��m=��C���O~��d��y��g�<��3IRu��F_�.�C���^�"���U��(�7� DP�<��8r�OXU�*M T�нl��+2�f�xr"hC�>:Yj���nC�y�!��qP���O*�	L�9��c�j8*��7����2'�o��_U�
�,�<�/7KJ��J��f��خy��f�6����zg�Ri��?4��#������B���S��{,�~��T���Y�l�׺N��Z��O:z�Ҡ��C<������I�
�v���k��=��$)�zuq��&�@9�x��ܮF����{p�
��#$R2�P���6F��3_J��=4�p\F:��~� �VI��'k׽_eq5�ͺW�ӧ�:a�%D�4�+���7��PL�$�Bėv����R�F��;�s��̈s=��c��a3�*rԆ�_�ʓ.����%��A��0�!J�g�ʾ�H�6ߟSJ���x��"�@�G^`F�����
�
�ZOc�> Jo�[tVZ�cBO�����l�ם:�'��GkN�;��O�aL��$��>�.�ᕆ3�����ȵQ�
|Y��e�,�{\��lޒ�rs�W�杬}��/V��\��łPf���6�����t��������C��*,���X��#x��!�eʊ:�ۊ.k���L��b�r��N���
����.>���t~�͵��׻��$b�L�[mzQ�k&G��emA�-r	�T�S����3�o2.��H�@� �A�[U�[?��8�(�TR�h{^o�$k�:�8z��G�Y6�
LɓS�>6��OdC��X�g ��U~��
!��"�g"7��%*ks`s���w�aP�31�P�����!RZ�ű*6�0�H<�3���?�{�X����|�)��kEO��G�l�
pϧN��7��n2�F�"m��e�����
2!H<��l(��U�����qÌ�s:]֗�c3�~2��B�[a\_�!�6��t�3��.�u��c䞹�T�u.|�S����ik�0l�!�V<,��-��k�|���=����k!V�E^팡<�U��n-gr���L1Lj��7��?��PYD/o�W"
����o�5���Ν�;�a
�
EX�N�Y�����VO����Boz��9��C���"���c�n�5bRJ�}�(�`��1m�%����߃�lZ��fC(P������,�.���8Y�X$�n1몚Ӟ��V�bc��`ec@M���}3ղ� ou,�<��E�e�a1��;`B��j���ms�55RbgC�p���0� �<v�z�oδU8�����ntyDs��L��H��?���-�,L?��G��u�ҮK+��zK�0M�VQ�B�){ϒ��ov9N��~<eyd}�"^>���"	׆!֊q�ʴ��]cVG��^�Y���B���8��#�H,�,��#��Q!n��ị�!�UڊA'��������<{��\�H]3�������?�������%~^��2KY{�w����;�i��^�П��gn6!��J�d�y�I�o+~�����T�}nO8��96�Y����gq��e��\������y����V��R�I��j���V/s�n1<=�$�.j�X�"U9��#Z��X:��(��K���r���:�d_xJSn� n��]#�ǅ��6'+��C�,�ly��ĜL(�kGcJ��|�;�H���}rcCX-��_����F�L�r|���o<v!����<��F�r��*��W�D�[��EH{*��2Y�K'���~��	{"�Ĥݮ�)Id����^��v�-�]���%0��EQ0s�X�����[�C�ՊM���T�S�?�(����������4J�-O�*�`����4����dȠ[���M4O'��0��XU����{�?�"C��v.�ݪ,����˛W.���4Ķ%�vXH� �4�FG
D�0<,��(p&޳E�E>-}� �x���	�BxC)�naet+}.�A�\�	Cc*�)�'\�]B�+��h��ӣ�-�Oӈ��y�j&�Jl��3b��٭�nP�T5��5z���.����VEϷ�E���=��"���%���%�3t��>�Z��G�k�|OF����=^�nh���hV�.��7W�zW^�5��y���=���f�2t��K�9Zl�CeΔ.+'�l6x�'����]r���9�9�	E�`:P�V0/k���$��(I�%e��t+���o<N����̃7'�L��F;���S6��w)
�7	�:������_ּO�R�ga��٪5\��������Kw��$@T��Vc�2��A.�_��I�J�g�̜|O�t��'�����?v	�q�8�� ?WyJ	H�|9����^%����	����[i�i������D�!�P*�#x�K�����Jz�����j��|���"gj� -�t$T�����r莨=k�w�H��y �X�������˔��,}`��*^�iV�$�3s���E�ݘh52.�]O�=�u��`�?,�|C&b4ݛd2*@~��6�
������G��%?'��Y��,4jQ��)�����pn��bu]z��^�e5���O�&��1��`f���J��@Z�h`v�$F�ۊB�;�n����2V@�3�3����؝C��*��Q��i�1�\��Xl5�o����.�]�V îL�S`3o�tW#���>=���T�d�޻fĮ�t�� �/�}:ug6:�,��u5w^��N_��f�R�흗&z~���~�ǂ��w�ҷ�-�Zu��nyU.��������9�l����ʢ8�p��,V��= b�۽�w��?��]�$���i]���5A�r�Fm�Qz���R{�:G.r�s�����^��%��t��B2���$�Xi�CFκ�ߦa]+cc�~�H�A�A�$��#w��3�(�V ����k�̪���i�(���"r���m����s!�P?JwM�}W�"^��M�ס�PZ�m����O��#f~樰���%�]��c�����dbn���?�KZ�`|@�ڃ�z�|�4;b�C���{�(0$GQ��b�g�UP�w��텤U������M����0���<�[��ZC�������I�cp3���t�aK��|�1i���w�1�='Y��总Ya�$���D26��5����$>��*㼧�QS��OP�	7uWe�4j�1��~��Z��M�?%�75� �������j:�TKia13D�V��@q��.�'�Vt��(fb��K�'�����K��{�TÛ$&�H�ֻ��ل����v}t<R�ݤ�8��Y��?�`	���`o![�������6Nn���&�y�fr���f�HT2�6q�̷A�k�"$��؋�]
��T�N~<�v����գ���<]�KT%0�e���,�lMr�����i7F#9�yn;�P�{bf^��;�r]��LaL����Up,�gk��e�b�rEqǼ�93�Eј�1'q%���٢�@��M��^����H����w����j���ec�ch�V�n!��\������\�?�9��d@���Y
В��	VR߸���i6�p�!h��j�q{�$1�]�>�\��'�0����5�Z
f�׈�o��o�%r��'�aFx���]��g]ʠ)����ܾ߶U��=�{���pywM��A��0��}\�`����vQ\�� EO^k{�
��iǽie��$�r��+z(��:���a%L�(p�f�#E��(S�-�7F�i�ߤ�@.�:���:�*����8R.jO��ZZ$���Sj���Ւb�}��e�#�,gQ��f��M���ʔ�����Fu8�o�wkk=���-:�v"��`y�v�b��nV>��c*�����R�_j�+�cz���#0���|1�oUV�t�6����J��0ۯ��{��Pj��9��%��{3 @����~Z	�VڛK1���>dF��[�I�0���'�1��wX98�Ϩ�WrB��d
���
�4A�?����~� �R�L�f5��7�j�Q/gu۞}�J�;��Ϗ�_	�&���魈�����#�z?a2��[�Y��z��F:�B�(�{
�G'���e']g�,�X�\�>�xl`���SB���㋏�!�8G��� ��%ɔ�c��� dF��_��hN�����n�sDdC:�1&	%?hضx�],����Ώ�Y:h�E�O�v.IV@F�#����k���6,"4=&��,ܓ��z��,��f�Vy&x��уx1�`"DId����L���*��+�1����LH�n���"�<}&�(c"}��� ⁲s퓎��s����9C��.{�䐚����y/7�d����6\i�U�+��0���[��K��f�}X�G�]����Vʀ�Z`Y��a�1-��9������� ejg����gm �N&59ٌ,g�����L�D����D�ο�����,p����&��6�H�����e�?����:��5 Hl:vTJ�>�]���2��J���C^�F��˴l��w�?/�s��sѲ���x,���ڳ��N�1@و�{���P�gf�w�1G��S�96r��wx}��,*Q��L��@�`{���>,5���M���)t�m�3靨���ugU��y�+A�Z'F��
�y9�MJC�JB�.}��%{M��Rd.�n��&3��[���Qڍ���>�!�Z����f���[+��	��qXߎ*MN��)�ع�	�3�\4E���b�X��V�[�1�֖��k�ku���*6%?����|ަ��R��ޛ�o�#� S�x���uB�J�I,��u�4������n��e����]���Tr��7��0�6�	֞yJ�N��d�;:3B�+n�aum#f�	G�lwK�	k���\��|^��#��
��¥R�+������Hu��G������gu��;)rƀ=|q���&&m��������Q��{`�J,C�!�ώ6����s!��.I{nCg��f/��^\�4l�3 ��h��(聹�h-1������&� 2�OӰD�T��������F<�)�0@�����K��K�<8��o��r�7�b�К�(|�D)h"���]��8������,��-��;�������޻Y+��QsN��%`xP���@�Ĳ���ʰ�����e�37@+q��?cN���:�O$��N�+�8o(�	SJ#��Qw��z�+pD�v)�_$��\-�ك���ۦ2(F��Yԧ�oי[�O$k,�2���0|��8�U�9�D��DtV�@�`�/QZ���VϦP�=	�hf�!}��"A�����e��(g&O/�j�F�v)�#�8�4j���~��,e<%���|����W�L�:֫ިp���iQnnD���i�Q>U����-����18����qȑO��&�­*��M���B��L5#�]XN�U ��������q��t�i������y���{��%ٝ�Nz�Vg�9��KJgg)�v�OS�mnC���(�ρ���]uD��&ͨ��0?Aj�������>����p`'���$d}��.V��{)�*�]�]A�� ��2S4�y�	�����,6����c�
��"1[`_�E��W.���-Q�R��M�,P�xx�}���&�qU�@Ñ���9+xJ��l��>
�%�3�����Co���y����<r�B��@��P�2�Y��S�;":p$�J|p�
�Ж�����ϵ^��-p�Q=�Hy���Qf9 ӭ7��z�V��52��zTV�_���Tݾ��F��h��l��=L�9Y��
\#�T���P��v�=�X<vBZ��Ց��e��y��%PYx�Ge���ݲc��A�4a�������b���VK�ƿP�d�/��*���Z#�KL0��1	YH���=�ʋ��L��f�g���.ނ�:d-�T)�hA䀐����A�l�Q�Lo��u�B�:�����i=C'Ba�)�ɍt���ٗ3%�Ծ"����ZG�sgBfM:Y���0O�l��H����m��Ye"oR%q,�K�7GI9♒^�P�[_I	F�#G�q5���=Kw�p;����K��\XWhݜ�'�ȸ�AX� ]��2:��{�r~����Q���U]�j�'�N��5�����H�l�1R{Ƒy�h~�ר�y�����g�{>6� \�,�P�����&���jך)=��˅%~$̏�i�O��s.(�`��T-��P��V�" ��(���Zn�;���"����Fe౺��)����dV��b�V2�q�6�l�#�{0�_�ہk�V�ջ4��$&;������,/���^cx�y�~���f���3<��|����m'|��Uw_ې�R)RE}�"܂���K��\��SY�~�j"�C��+�($g�:�ښ9Y(�$�&���Y�6��@�ՈD���r#m�q�;C��I��� �>}RuĒ5�$��I�;�@q-�&�>��Le��gr6@���
XD*���ƭ��;��K����y�"c�5���}즂36����FA�W?�[;��C�����e���0�a���%_���UިMw~��uj�p����"�x�-�C�i����'�L�GWq
~��anf�%/<z04¤+kf\ȱ���X��^^��q)�C�9���f�ԕ�+�X����c����~�O��[ؗǦ%�Xj)���s{����"=9aF�=�o���u|1&�q��%W1ʚyJh8�]�T�"ׄ~��8�+:�˔��i	F\�Wi�ЗGp��8���I���H!��Ƴpt6�������}��F��T��