XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��|
{�\ J1;*�E�C�~?��;��1�³���$.0FȾ�}?~�����klC-��1���۝*��Gs#��R>���p�x�YB�#IO�^ RN?;K�F���6�_�A�w��x �@U�3�l�R�+�6�����`���T��%��b��H�E5a�b�-�f^����%f�7�o�l2S#8�RQ`�@8����1�X�b��-�c�*΢�Gno�FL��u-W���3�$`p_;^�{���«W��ʿ=��R����1P�(s��7S�-?������a<�mӋP�ia��������nML��l>��+rb廰[[g>�u
��p �₂�Dy��ݍ���	6�o��m���6���#:k�Ȣ>��"p<�}���r�_��T7�7SEO�I�|҅o@H�lYW��p*t�|^�a�ϧ���w(����H�)0��R�5�(?���A�� ��7�T�˄���'y����+v/bPmپ�wg��F`6a���\�mH�H����;����ley�k �N˦45��5$���W�p�w��#��Q�_�m�E�9��`��S�1�?��
,�� P����JE]7�J"q^ ́w��_5!	>HG��9�����Ӫ�2��!E���`$����J�Q*~\����5���4�ݾ�w����T�pA;��3�(��$� �1p�cd�D�۟�,&v)�l�&��s�z��^F���wɩ�~�����p�\��h��$��a�8�淳�o܌���N��*A5H(���=XlxVHYEB    290e     af0�pΦ�Z	���=����*	�J���
��?6wq����.��~�3�M��If��$!������4+�$�w�Qn������/�\��c�o�$vr�l$�|u1ˇ�_���Z<_wKwP���]+'C��ћk�Hf/7H�qZ幛Yz��5!�ш]�7�Ad�)��d��m���D�A��r��X*���w�n���Ȁ��*Hp�cs�E	�w/�M��\4�(��y��C'�FV?��(�(��R(�m>��e.�������յ����d��G�.�譃��i٫�=�}T�9Q����<
�F?�du� �"����2��*�ЌdC����W��ECp(�͚b���z�a��8�Y�R��y�Ξ�|����,(.?]-I�����U�P8�BFy����Cv��ٳ����c�_�
UA�Rqe���s_h��=�O��F��9t��Oʷ��o�n=��5�t~���a��+5=,��:���n���{c9����hTa�2�7��wC��g$�r�fzR�{O,
��� R،͌����(连1�6idh� �@�`'} ��D��[' b^��*�GZ�4�Υ�5a4-�I�$j|:ؙKAF�bh�8 ����Q-��(y���-���~%9μ�
>����V_GcqA����0L��/�\���I���ZZmB�9�+�)�fe��$D�Y�� ��^"X�6p��X��6QJ�ٟ�hӎ���&�Û,;�ܤ![���U�`��G���uP����'�P�Z����O�U����[B�z�H����QaI~��>��NcY4dA��đ��7�kd�(X���X����;%��)WZ9oHoD�>�$��LM����dsw��y&��U��t�Co��'�LL�o Q��ᴄ �wM�:�~��SxX��(ؔcqÐ���N���s�C����Q,�B�MЄ��ҭ_ x��^��!d�����x��˿�u�Ⱥ Ϝp�&���+q��)��]g-u኶��"`�H�Ĳ���H0�����	�r6;�����_	� s1��Lȕ��W9$ֲ߭��Eι�o�RE�K�����L~!A �N�������Y:�7BkRe�T���D+8hH:��bC��3�5����_W0� ƏH�"����|:}��J.�\hj����G6"�%�.��B�h~}y>��_�:���|BLSQ��)Eֺ-�J�v�עqv�O�Yt�q����c��4�GY�%�Gi_�p��A�*e�ݬ2 ��h�o��q���l�Q,��uD~��3����d�
�dC����x%T�q�G�0���=qr��*M��	}Z�b���Bȍg'��0Fs���.�"�����-���������kOOc٤���<�y4 ny���+&r�)�y\`$]~���@�j��e�)-�#��*��|��w.��/p�h�^�V�	Z�V�]��PQ�V����m�$]�<��t@_v�D�b8�7��2�k`�
���/Z�x"� �L�J��KB�0V�a��Г��`"�F�>����8��"I��W�����͇�A��|3�s?�J4�+��,?�F_X_�(�&�sK0lww(v�ˣ}�ULse�-�z
l����-=RT�Mn�Ԗ���?M���kOyF���\�>��=��Ѣ�q˫n-���K�F�N���F���ʂ�<��.V^� �e����>!� �� z���'���Jjz�G�������F�2�Q�7��l�`�$��t�⨄2����]�2�R>�L�5N�ǎ�����ʩ�SS�~s[H"�*E6Lū�V5��d�S}��j�9�D���u^I�ފ��x���l�#�,�[�^N�����ж�NM �@f��s�R/&�;���$��7};y����x9��x�0�d��Ng/:����m�Hm�5.�d3V�T�$�$ϡ�w/ڑ�-��e�T{7?:�)s�Ҏ�N2��1�齙^�/[��,{"ԧ�+'W�z�+/�l�+~Ҧ���3?i�^�
���Ck�����HJr�5��'�̥Qaq&��L# ��l���E�AK,�0��( ���Q:P�oK�[Nr�D�c�G�/����1�uԧ���
�0��0;��֧Nw�!'�(�X�&ܢ�ʸ�%�(>��$�`"���H'
V
ª_�;����B����R��|N��ɧ3.��Ʒt�=r�\{�l��Y�Gߴ�Hk�޺����*��W��Lݮ}i�kȠb�d�j�ЇJ
�w��F���7 ���@�q��iQz�����Y6��R��'�.��[~�=P[l~G޴�'=��rM&�^i��[�<Q����a�`�u��?��JC�]���Q�����k6˃9���J%}7�Al��ؤ9�E�M�J�g�
~x�
��a�m�Z����ގ�N��v'`�UtrE���F'�ףO��ϩ����x�H/$��lCyI~a3���ew�#�7Nl\R�Fae��B��9��K�u3-79����[g-�~�;h��Al�O���㚆�v���ΰ�u`0Z��7O��	�G÷�K�>�h��"1��I�=�c����5���Anno��(�%��V�0�?�K�yК���w�E��H���jdz�Kp�K�y��Ss�)���<�g�Ĥf=�Ap�,c���)y4{༰�p՞?P�Ᏽ;�7<���#I:�_f7QԽ�� �ꎑ���A���X'7M�F�N$��ʙ5N�WM���1Ŗ��JRj�F�rHӆT� 1yZO0�!vǅC'��Q�P�̊+�tf�