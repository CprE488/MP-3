XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��L�VV��w�:%��(N5o�at���KX	�[b9n��У	n��&��8�ueO-���w�p)�h{ȒJz�uV9�8��"�o��K/�K�kO�']2L������B���y"򳩸ӾT��r�a9�5���~��0)�`��`�2�!o�[������K��C�C���wؖ�#��l"‴g��$0�{=Й���3��|��lwSt��ʬ"Ӿ�g�����{-��<w��uE�]a�1�!�+ոO�^!�ԤJ2�y�Մ�u�J�x�5�:��o���߁�������C-��avõ7V	 �y͜,[$�T�`qC�>|b���fOW�`��L(�/�ܫ�ɴ���`�u�I�8�D��JmduL]�5�թ������Τu�&mk�QH�6�S����1�f��ѳs{^���{D(K�*O'[�\6��NKZ�<r&���7w�A�*��
[_�M}&k��fT�i��3�;��Ĵ[`�46�}�p5u	b[��Q(�SK)��/�3���u4�R3��'3��j&�7E��P��������7
Z��"�c�@�c���X�\�R��vp�-ŋ����z�E�#L��L�� ��9*Ж�_y@�T�ow�O�}m�ά:j���2h�:�LuvW�ٍ��r�p��Bn�)��Bĭh��-m'ti`���|4�������2�(yL2i��{�C>45l��ʜR�j�?�8�����8��ϥSP��'u�8�[��qF��V�ŽN�����J��Is�0��Lw<XlxVHYEB    3a46    1050�����&��;���/��舅��Y�6ڬ�w`�U�N�S�at��8���rM������QQn���זh����~��}�+K'�>�V�!��h`\w_��Q�OjmQ�!�Wqk�f"���(��}�T�[�ף����Fx5�3�U�KΡY�[,<�1��9ʽkQ�$���t������h�6*R�>8��'��>��i��a�^�V�l s���u����Q���l�RT
����_lw��Q����T��fg��Сp�����?�
����w��O�����`a�}�����mDK��	��I/�N��H핮R��H��{I`s��I��q8WO���Gxֳ�K��P������5�i1z�c-�e"0�AJ4,A?��n�(�ƙ�f�N]I�b� sE�]X?/�U�񞇼��Ufw $�Ɗ���I�̛.pi_��(B�>��BHm�P��h%��LZ��F6!%�i�&g�x���H��FY��M�	"U�#�]�,��U�Ja�;��m ���W�Se�����A �_YWһ�r;=�A��m��'R���	0d�K]r�8y@�	�R�	�G�g}1Yd����!�7����������������K�{��{���5{�,Da�X+^a❛nk�5#���k� ��>�c����hݭ�E"Lkc�髉>�Y�}	|"m���Q�ߥ�_G6@/�3?5�eS�GY9�Uwoe{����}?ݑ�oV�rI���x��WQ�&E��$na�fw��b6�z���h��x+��p֟����nP���	^���\X�\-��=��Yw[Xj�!�ʋ/�4X��E�Ď��{��N�ǩ^zv�2�Js���{}N<>�m�W��@/Z.$��Ɵ�]��}�\�wL;�3�0M�rV��=�v�=QM�vJח���9��;��'��x�}o=����T�ůL�0o��V�b
$_g�dܧ�	vq���K���������!����{8��`R%�� �o�x/����1#�4Iq�`�X�oc�.�����{M)��,�����4��ơ��4���(6���{������G`}4^Q����*���"����Bp�?P,�AS�F'q��H��"Ȃ����|`D�IJ�����_��_�R@e���q6��k_ߪA�=�tn��8�8�<�h���=�T�^�N8V��|�Y@�D�si���T�KX��|�ESȶ-q�(�]=
̊1��jT����׫NC83�a���h4s�}:�rN���<�ӌ#s���ۘ��e��%���#d�"�3�d�w	��AqclXC��ֿ.z����l��K��{���W�"�g6]��5H�),�EE�ߺU��oD�Y%��"M�>�!����@x�I�!1ϳ�W�E���x��������a�]ѡ�N�Ь����&�A�?��LU��+x����L{�Ph��?�敺P��tL��2�ǟ��e���B��V�/�z��1��� �ڠ~�aӪ�$f���T��+h�qZ�K�Y�|��'�KP�poS��G���_l��$���\�Oǋ}���38�C 荸UW�W�&�ۥ�����H�ܥ�]������aй/����_�K�h�qk�ؙ}���J"�Rn�^05�Xd�TC��!�='�p	k��
�`�ҫϠ~��d���**'����z�3R���A��ƮV�Y�*ҁ.H��3��J�*%�pi�~���0≂���k�s9΋j}~9�_=�l�?\��T6G�6&Aw\d	1p
��PY1�>	�����=ߣT�Խ��@�������Q�G[3�*y�C�鍦�V6�zo�H?@��x�e��r�SK�ab��UUU�#��/Jo�lT��O��re�J~�fS>ˑ6�"�Ń�5�_�EhtІ�Q
��ص)���b�*��ڐ����%	pT�	���h�aOD@�T��]}g�f3�a[�r�>��(��g�����드x���ü�![�:�t��N���gHV���ɽ��SP}]�`��Ɏ;
�����C��7�Y��{
K���huF%�N'�2���P�yƬ�D�er*P��U�詤�#��<^�$ J��ZhL�"0^���Q�RI
g�D����!fb �=�f��� D��W?o�(:��==���0�}6�եyt�� ����З��X���Amw_2���>o�nSn5��a���+lea��5����u^��ȁ��o��f���َ��I��q{�%�)�$�#����"%)�]$�! `�Z�`��_�L��&�×b�w�x3Mc&������G���}�6G״��pN�#�>���~&�����,�	 ��7i<��eҎ��	��3AB*�C���݃�z';ؖ(wϾ
����E�"هp����i���{A��s��
,)���P��Vt�Fh(fMv�8a�xi�����zcNSgマ�n�;���
��R�5��}�X��|��4�8X���]�Mϰs���Y����۪ VO��[��{,30}�U��A��M!]I=�|r���v�4����U.Y�T�y���]�@[{L!ЉJ+�:��^�����)YW:���,.`��)>dv�����PD���.��hN�]ب_��Z��/�#��	�ܼ;&��R�f�'IO���B"�$>cY�+�/ϱ$���H=�3!-����$����6h0I�/�>�hX�;���f@p��O�����g>�B���j���hX��I����Y�b4��\�����>�7���|,��a؉���*x�=ð�P�g�Z+Q8�vx��5:]H^Tiջz��2m��*v;��M<�1*Skz�^��I�o�Ѿ[�x?���l�ף	z���ǣ��]>M:w0�`�m"�"��U��P���-A�[�����r4}1�o�SH3)4fSb��E|^3m�/�3�{U�lX�(���r�Ɓ�xlWŴ�OU���ʜݢ��V e4K�\�����IuuC�UB�|6�KH���΀��eeY�G�<�[?GA��s�gF��B��m����Gg.���=J�&r�GC���Ҫ }�;� �fb�[;�<������AU{�����c�M'т����p��8:?ǲu��i��e���0��A_-���AF�`�
�}u�e`a��(+�͛.6��<�3�lm�_E�j�ɿ]}^��3�dU�}:��=�Y$@�gtm�"J�^����j���wU��ZO �.�YUwF
�e��£�
j.���#�CTg_����g�����U��㆔���/��4�	���	;�l���[���,�mIJ�3���{���ϕ�ݍ�q�fkP�V5:e�������fDt�3�д��8�;k�E�3����I@���q.�oyAQ ����������cG3���d�V���MTz��ӷ2�-���4�40"^$~�C���ҟ�u:����Ԡ�J����zq���F�n��<�qr	�I��n��	�b�0�dK�V8w=k}��~��Y[␌�>	�Kt0˥�`[�Q<������ ������Z�ܻ�Qԓ�:��V��38?��k��,կ�7T��D��Y��~H���R��7�:Xx}�X���2��B���M��S}�4	��	��)'�����~��Ҁ"�.��lA	�8�a'�g>�M�Νpj��#��3.��������L�\L��)����`�>�փ��nކ�A8r�q}-�[bJ�������W���k�H�w�
!9�]cc�ЃH�aНn��� >hY�Wʫ��D�s��d�rY9����ͅ����]ԡ�}��ӣ�%�<�k�`���%�Q��!���?�$�Z1��Pv)�f.E:��B���+�3���CX������8,+�t�ٷ������	�^���e�G���.�$[d'2�T�<��c��/Mug2�y�k�3e�,,Ƞ0�L��&���A
��*:9E_��6�n�V�h*@4,����?^H�M����KaH�bX�6�=j���N�Y7r��$P�u��{��,�z�^ۯ�r��2����Ÿ�Л|˶B��S���Ц������?�i/� I����n� �O�>�G�ѰX��=1��=��VD'#��m�E���4w�j]��_�!���K�