XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W֏��񼇘���4��U몺"�/��RX��v�	v����$�6����ţ�m
��s.^x1��}pI	���.��A-�}P�� ����� �!�dۙ'T���+ĄĚ���T��+�@�$nb�j@|ս_��6a#?�Vʐ����E�i��9�R�t�o G���
*�+�����a�R�m>P�ܳ���L��`��0�.��\$���=�a��($��áa�DU7$��K:�_��$`%w�3���ҷ���ڹ������V�E,��3+!~����[��S0���@(��SC����1�9���E"����R�}+���-�{�?�N�;�rk8aJ2�/��]�'��T7q�Divc�t��B��r�e#����G)F�� s(Jp���?m����ǶS$���<@���U�y����b�Lщ��+b�Q�؀}qP<�H�Fr�03�_�9��@������ݯ�����kZ�u�κ��|�=
�S 
D�D��5ͨӀ��낲Ii�/��>m{��3&yr���� ТM�;�	$�]�;�.��Q.W��rߍ�;�lK�c�%9m����T�?W�phS�(\DY�Ŏ���!���T�{I&x����7���r?��I�;_�������*|)�k�!����-��A�ONq�+:,Nuz\��B	z#50`�Y?6�7����_c�%3�p�e*��v�(F�����+MآCO	?�v��D�`�\w<��`�ڬ���`�M�DX���pXlxVHYEB     f9d     6c0�Pϔ�)���/��p��U<�Zї�A�j/�k�1���}�%& ���h�Dx������X�� 8���s�4؞�S�k�ƥ֏8�0����(i,��.sy~���P�qԹ?&�Y�	�_�(ɭLN�>	3~]�� ��!2���Gd���1�\uBE_�q�6�J�(�Ӹ-B�:z�P��C#'�vy��M'E�%�R�!>^�D��F��
ᵅ�uף�:i��(9F�h�T��be�
i�@�6�Eu�M&�{��'O*-��\��􃳷�u��	ۍ �������g�G����!' 9Ϳ��������K���ΉX2�������m'N9ĭ�ꄄ��k2�1�>�6�M'�x�ی�o|\��Yh����lg���� ��\	�Cv��|��F���e�pom�P���n�$��_2�cS!+���k����D`�zv����6�p�� ��n<=���
~��� &��ǎ�*����ٕ��X�j�1+��`��0j�b����F��u�y�k!�5�b'7���`�"~r ���(��Aſ�o�9�gJ�����u�k&�l��N�U,�]={fkٕ�>#�ڶz�+�˫lt�� P3uH�Kc/X�mw� U�Ug�C�t��hC��'P���ZC��J���ǐ��Xa��*uV�:tcK�ȉ��.^x�9�eTV8�����M�����6-�[��,��4�c�����=y/C;9�?u���ZB#�a��8��)�D~�le���5���i�n2�nFH�>�����KB�~�.��m�Lf|���)gGl��;��2\C�
�v��;�y�w�T0�n�t �;I�n�?�B��a�5c�hY��e�ޠҬ����6d�j�K�h�١O��b�^���+��ZQ}b���w�`j}�C׸e�H�
ۼ� ��ί��Sl8ڨ���W}�M!�����/"f8qTkǢ���v�o�h����-}���Q�H�.�{�➂W(�d򼅅�Iy�Ύ�X@�[/���ko�4"�է�n��5���^�b"�({���
��]�kV�\9M��wco�*N�ʶwŽ9��\+`T3�e�Ξ��!]�G��5�f�A��oi���;,��##�L��><kwi��3����5\F���Ą{�j�ڠץ���ć���r����kT�z�2�{aE�t��:a�2I��l~�*��z_�����p_��s�v��=3*�n�ɣ$�<-���+ѧx���Il ���*�Ts�!}ǩ{�	ew��_��;t]RTH���G׹�����Ø+I��t(������'�8N��C�ê�Z;O���5��X�"����~֦Z�U)?ڮRi� P�{-{3	+����(9�F��٧���#z�QWCY=��Q�-ڼ�LPB����
Ǌ��\j��*"]�,צɀ$P^b�[I��û��L�C��� In��7�Ƀs�P�w�7͝��q�llP��6��g�8�bxӿ��`R[)��(�4W�^��S�㩨�)��87����F�k�����_IR�BWC�Me��"�x�qN�6��p}�E��D8�LʽӜ}�E�y �+�Ċ�{����終�m��?�*'����H%��B5XNR�z9f�����O� �����;e��Ȁ>�-X����=��"�&{o �SN��6��sQ?Q`!.{K���rQ�D�!��җu�6d]ѭH#�