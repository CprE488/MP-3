XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����U7�}�E�y=r�x��Z���̝D�G�O�S����f�7?G���y06e�I3e�U!&`we�?������S��uWHt�f�8:ˍ�Pu)k�����V�2u.W�;F�t�X�}���c������
��,j�^���-�r\���/�e�9�Jh���oĖz+�S'hat��oN�5m��_����7[���7{K.�Z�ϥ�|�8�	+�?��Ր7��t���+� �x��W?^���fV��bKs�D!z�B?�=g5�DG$���N �(��/����'U��ͭ������w��0r����/�aR�;4~6�B�\�֮��CT�U��rSU�3�k���N������;���ӷxJ��.�8�J����ʸ�v�ۋ8X�:��L-�4?�~�0�������=,���c�H	��}}����3��p�z��G���u�,>�t�����ƀL��Nq�̹ѰE��Y1,�C��I�-+���;0(bӭ����h&��.[���z�w�Z;�{�uf�&����c?����_h{���i��9��(��% /6�{��eMѐb<�rA&���,xrQ<��Z�m��>��_�E�$�/�����]��5T�!�����z�������4W���O�.͘4ӎ=[�Ѳj!�yЏ����dusM�z�^�MF�F[�ڞ�A���a$�e�����A9��w��}0��Up���;G���h⺶�?����T���YX����@�
7YXlxVHYEB    82c3    1970�Z��lnn� ,{-�fu�0�F��x�C�B�;��|�^���'��͠z�,�����~���i���6��g�ǯ�����щ�Sŭ���T�rYk�~w@�PӲ!5RCp8�S�l]k�C����sS͗-�L���ZU�$DS��ܝ�=v��:/g���w�]�d0�u=�=�I ��V(�]���{iW�|;���$ـ/�"d�(E�V4��9���vAh�/
���-B�MF���5��b.~5���@k
O/�� Bi=e���� ���if�z{��D���bz�\�����>��<|i��AU�Zo�Y+�'qgN��+��A�4o�Z��1�&�+'̷� �Ƚ�tp_�a��?��V���ێR��&���P;/�{��g��v��(�fl#��� ��Z5L�vk�I?��#-�@��6���H��ĸ-)����L�(�Nu�����<��������H���d�Ȇ.��#����� ����mzsrWK�� �S<{�����p�H����{���t�a�����p���P�AI�{��9o_��I�v�����՚o�{�Z��Kpu���s(��TvO�%	�>�Sޜ�r �x*����P����3� �Y,T�F�`BιZ[��AJ��w]����.�x�)�����(N�y�>u��s>խ�>o�z��u�S���G�$�g��V����x��j/x�9Y�(�^h�CB��<a���U�Xo�7�s$s.1@���C/�8�\'���E��(��:��G���ѳd�.�x���:�:�����M,����|�\��T�+�qI'���n�����U�J@)co)��+1��%�k>�B3��r�A��$"׻�P������\��/�{���k�"U>��� ?gg��=|�������v���v�,�W�R��m>!��"���;��oK�Hr_�9��q�$�s|�e�mV�e�O1�%�z�Aݶxw��=ک���e j'u�^D��H�ꨲ9�][�F��cZ��`FZ�"�(.��A����`�ek����c��3��I�w���(����d2����Ɛ^2̳ l���>�l�OU�SBi1�q���|��$`�Wɫz)�{�6a�<QP�A�^w���ⱄw�9]g�ܘX�g#��:z����p�{�H�㨑�5)0d�I��������;��Х�$&2�Pg��t�T�/#,�(lԘ�)K-�W'h�n�,C�T)�r�X^� �@1�O�܎�2��GuT&\s/�}ƀ�����^�m\}Ctu)%:��9v�|9�:)���2��n��b�Ɂ��EA�"�?�� _ 	GD��s��O9�M�����$8�ng����Y-(��Z\,���Nb��.��D���_8�Ħk��G�H���q��V��^{��op~��p]�i���&�@1��;��9%⺈p}��Br���̿iK�h4�=�-̡{�T��?��瘿5Z?�h/O�C������M��o�4�܍�KT��! d}kV�mq:'P���l[�j����*�a�����A�ؒ&�n(�-��ˆȐ�l
�go-��d�w@� uĩ+�馊~'糭eC�c���e������M~oL�q��/���E��I]J�yeG�U���"�/Q�
�����V�$���{��'+��S��f�Ѫ�2�(��S���;F\��L�L����J�Z�늏��ѕ��C���m���A*���`���iR����k��=�i�����F�� mvr�΃d�`��ЁϤc�\�4b���"��Q=�2�:&�Jf�/�!�}@�fO��f���>�i�A�%T*989!��0���F�kbx�I>�����=�4��  �k<��?��ŏ̈́���1�[�k2�.]���ڠ"����ƓyX[UڔR ����x��tTn��v�8�Vς�8�ul}Kꬡ�(�����{���#2��a��uD�Qv�8��H=�L����/W�Z�D6��V�rJ�=*+��<�>T�I5[!��"�����"#NX�G�	���;�R�� ܸ��&���k�j���m�
 ��[8=s��b륎��6�|&~8��5�C$q2�h��4�ǖ�!HP'љQQ�5YN2F�Q���Db��)��M�K7������)�Ռ�"QU�b��`)	�J\9��+��2��D�-PЈ~2�9�C��77��Pv��ʲ󅥐��q�r�����q�J��X^sK�$6���@���k������6t�kʸ��N."ne?�
IAxsGج���ю�S���Eue4z\�u�L�⎘��%���� �a��;��љ�l��!�W��L�^������D�8�r��c"g��>���u���:�п�	Ub<����� rEAX3��bG�e�2���x����Q?÷�3�ႈ��n�ɷ>�G7��9��S��$W������1��̛�������ק��̮�m�ra@�ϻ8���"�P&C������H8�L�ɑ��Ǜ�S�d,I����}+�Ǥ8J��lK�z�K�b��g�ύj�M�@�<w\���tLX-K�8LL��Ύ���U�KP�<N��)�f��۵�2
��A���)&���;��t4�--ȐU�TdÄ"8��gˊġ�@az%_<����|b'-ԇf�طoUq�E���L1V+|-�˕r��4�~	g�?�CS10u����"j(�n�"jE�$S������k��0��Sx�&I������AS%詾�/+å�E{�� �[ ��{�uغ���������w�YT�n�қ|�X��8�L@��j��B�!�n���uZ9��za7D!؁P��}20ݿ廍h�������z��3�E#��'���+�ǯ��׼ M��V�|�蛙���/P|BM���C#����t�K�@%�%|0�)R�7Q�f#�fs�}�D��saj�V����d�U�-#%���=� T���#�٬Ka��
j��� M0@��~����z*�����Va��*.;ы�%�d�lY7E�S�I�;��vs�^z>��1X�-:-2��>�O@@�̷�]' �f�F	���_��\�oPRe~H�:Y���m3�@�ş���2l�лÀ�0��u�zm��J��R !��5=����D�Me.H����߫jn�hoC�Ygm���˨�0Gz7T���6��?�!G�;.ߕ�ck��K%0��Þc\�*�3����z	��l9����VT�y0��yً�wdp�Cc�k���x�1��������s<�\�X s�d����m���hqk�̛�		��u�ēJ����g�}X������B� ����i�R=;cq{:Q�0��Dx8���L��o�W���f)x��,�p�Õ�yN����L3|��@��$8/�v䝿Ht6"ۍU)8'��]HO�[�1��H9�"��$�v�|n9�F8{��ջ򼢨^��_���m�&��N��/E��;Sؒ���݈��5�#���]*�q���	�q��2?��,�8��e�vӰ�[o0�N��g��ר�W0��{iм�C&���&��~g$��Wwg@?�29�9�B� G�l'���{�
�6�	�e�"Q��`��2u/1���1^/�u�D�Nz�c2�^�	�|�v����<$���Lq���Q�*T�t�!9^_��"v��`8	�M	�2�f�8��餇�,�D�ơE]"����UHX:l �N���&ҷ�{_�М�	�CI[#p�Z�E���V�D...$�X��c�� %���f�.L*浔t��e����Hi����z�����Y�׃��?Op�(�L�ֲ����	��p�T�6|�J���q��- �νg�'�ײ�jX���DT�q�9H�_�%���f@��?���G�ʢ\<����+_�\���	9ӌNٶ��	f#���ۤ�l����8�
�䨯4tXW�pq�^(:RQ8�o@��2�΁���x0�
�QX8����$}��s�A���kq!��<	������\'�*���B1r=W !ۄ7Ď/kKes�W�y>����;@�ʴ`U�Z&��A^^�D�fM	����Z�(3��<�$'�z�ӕc�HY�lW�B�J���7� p�L�G�s#�����L2�Ĝ���,s�<#��X+�C�����$	��f�ܹ�T�ݹ���轂�� �g��)6��F󮁖T剒��/��$�;�[a5�*�w�N˒�Wt��R"3L���->�m�3�+	�"��&�r������"�����,[�M}�P��9��+<v���t��&�Z�C�e�w�A��h���$Y��m��= #�W�٣\�AڊL+�6��F�AO�5v����NlC���t���"��\詍�܏Mc�;.�(y�z.�W{>�A,+[Ƭb<�8,�{�/��l?�W�.0�esxM5U�)/�؛��0@5���|x�k�A՝(W��蠟f��4|>�H6�h	��y7���旞��)��=�.^=�#�[��ר&n�g��zp��^a�Y�4�1���}�����n�	&�T~��7��Z�|@���������<���ꛑ�2ABwh{\3�˘���)%�Sm���&�e��o��܎�!�j�=��L77���1�|��r��}9j��{�(����SU�M�w��mʐ�@�&��A���ms'��3PA,*����h���� ����n�I]1��d�Ǽ�V�	
�{����*�1���@a����!|p�E�&���a��.&ZB��7!�E�[a��(3�2o5�8����՛7�!������4���O2D
M���oڢ���J��0�uF ��	GN=�ϳg4\`��x��쳭�S{��O4�<��w�o�� �b��v�r[����1BAl���8�-,�%�T�����Qz�ú�^?�W�Un�[� ����ԡC�Ⱉ��h.���lAm�Dי��&��T�֤��:�9�t����B��-ߊ��G�F��~bg!HW����j��w�g+y�:寏 ̟<�ϴN��p �����U"Nq5ו������_Ʉ�0|���5e�
���'i��zk���`�,����@�1[-�C�P�,�I���'xE�	;~&��ǻ��CA>���e���Ka�������Q���hB潞�mde,�������¢����b�c��cAЪ { ��������
�{�P��*s0L	�1ʮ.]��ե�<T^�htCK���(>�~�*&1b�'��L����rͷ�Z�tS�K�XCCl��@u�Sd.�H�\�?xH�P>	`���)�3 kؙ��$�x}�\O��*�-���Gr7!Վ>�t�WKVU�+9��{�����/�����(����^ts�"V�z�����\�#*� V7�=f��t�yP��}��h@�+U��GiV�e�1]�G��s7��e-m�lޝ�#��+�1�K�H���ĝT/����$���\��3KQ�ܚA����������^��[��C�B��+Σ�]C��Y&JYE!猎������MD5�D!���e�8V�W�����.�g����֙(�����M1�M���8�F��@D�Հw$�[��<��$��s1}!~�l�و��#]�g�ݾ{	��'����+h���p��2��[ׁ(���Z+
f 6~��ᓚ��Ɂ>��T�YI�:�J��gL�Ք��|�2t�����ˬ����}r�%�,���~��@,��|�u#Z�0qd;��tq\~ɮ�yav��׉%�|�CE&��PѹL2����n��Z����9w!�u�g��8��ٶ[?�K�6�f����[#~�Ӽ(P�!}�1"��/�E�kF�V֋����7�;9sO-֘�H�F�re$2ݡM�B� Q�ܻ��	�D�	G2�6s;�k�`�Yw�a"i7��h��x�PP��� �V�R6��3-�<z�ZfĨ��\^VH<BH�aZ�����`y�N$=�[�YȊjWs��	���Zk|Jw�d͕߀yyg R!S�y[�I�{�DG��kෂ�	����A��V�?�(�M��@|o�ې2ۢKX�Qs!	��_~4�'+�(����	¦mT�$��g��	��6�ϲ�C�����<���%'�Ɣ3ȅ_�R%E�����LY�{�;F�࿵�sM ���SQ��`�����^�Y6.��x���X���+Vj؈{���>C���D;Xws��x�y�8?�h��yPi*b��)4_��H�ݬ@ሦ��~^�x#c-�"����&=�/ii@��?̞�B��[A3M�rP\��&�Փ��Sj?w�4�}=a^L��L�q1S ��>���d\���. ]C\kL,Z��+��wݓ��H�
�.�$7x;��`���