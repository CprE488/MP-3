XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G��2�ea�9AY��i�A�E�׵�X����*:o�+Q>i
Ќ�Ȉ%G%�J�ke�$��+bN[N3Z3�� ��x���}!�<�{gd�!HYS�s����N���jݥ_OW_��lJ!q�������_#y-?'�j�eZl�	Za�{�6�NW�*�L�\�ѥj�?b�.�H��%��c9Z����ч���ܜM���XoGsƸ�M2���Q}7R��Ō��a�t�;l	�I4l����)o�d�SD��+9]Q���_-�6V�iL"��/3�E���/r+sr�j�,#�=H6&�a�
嘘�f�u��H��Z��E/����v��*���)��__��:)gcSbs<�PRP��'v���Y��e�����1r����C���c	6�}�9�G�u)��h��b � �U�)����x��6�9]g�EF�1_4zU+����޻��n��e]a":t'��[A��ph�V����D�)��P�x
�P�5���S���_�%�޾��f��YL��.L�O$d>�-�uu5|�0�J���6T��c{q?���+9��c��H�y�P'�\�u�!��/3�p��z�O�ɵFi>��Ej��)���֊��K>�iz~��P�f�?mDa���
�O�_{�)F/R���D/�����'�sS��\����y���ZT=�{*��a�7��`��&�Y�]��8%�;]���Cx�g��(X�(���x �yKh~��n�����U� A�֜NS��XlxVHYEB    5cad     f00ѻVT����[�3R��]qm�;�"�� �]nR��[��5�d}Sv���蟇 V��.�o۟k�ล��yZT,��� | [lYR_��5�C~H4Gh�V�����}�s���c�n����V2���
��8��p��7�5s�V�:܇1"��uŹ`�#~�|󶄼�$�q�L(���J'6.�t:�8�?�ִf�0u}[���%�@Rk'�*
�;p�>���W��ߓaC�`sV��#r����a������!��&w ����E�6m}��g�L.�W���~��G�:L�9����ؿ��ZL - 1��J���!`�r��Z�J)n��H��@��H�W=�3����-m�z\PĴ�.������VO�#�����G$��Z�1��:�Ϟ�T)lo��9���S���93�h7WD�i���pC�� �^b����l��*ь��j������d�G)۔.W��Y�V�\�$6�ǂ)3��� :T�M� %�������� �[�v�����aJ��m�<j�Kk���
�^l�|�*.��I�sH�C)��>���4�U/�
Yŗ���i�BT��b�S��/FK �H �d;�F�9'��M_��$�E�`B����b�����46� 66�W����z!���_l������{0�5@&�9��*f���K�}	���R�=)�n�dބX��ha����Z�5"\���-�0"� >�Rw���Y�������aesFy���Q뎔���+2m���4m3�>��/)
���DLQ�Y�\5���@D�ffE0Jɦ҆\_.yJ�ܽ�^#z�y�&�B�r�,�h��h&����G
�ț5���� �XTs6�'������.W?�IlY񂊉�!3�$��¶�����f����݆HIO&3��v=<��n��63�v����0�y΁Zs"�ϗםLHȮ�'Xs2���l�Wwx�����N(�ME`6-��N����?�5"+-���|L��t����3I����D~��C�{Ӽ�Y�?90���{���G�A ��Ӄ>��1;ȭs6��TY"A��lx<H�N�g�&E8`�Ic<B5W/����u�kU%RN� m� N��W��XU�w���W����C�`�<����,���р��z+�j̑\�4��T����%����&8"|����M��Ԥ7tR�����0� ���o+����C��m�@���!��A�o�>�+]"bd�x�Y�s1��$q<iM�F5���.��,-�� N���<� ��G����
=mi9^��'��	2x}�'X�[��)!8�w[<�&{�ρ�gxnI'7�(n#�ق�W�M*�r�ч�t?��#�g����_M4AE�;�L��SxNF]�;'��ĭ��z0����b��Q����>�����WmqPG��tG�)����(3w!*.|���EaB$h[���r��ȳ〗E�8V�8c0)@��1��2�ψ�9Z�Ws� D,�ի<�:_#MM�$H�8�de�� �|����P��}R|�0s��N��l��%���ڦ��h���hA�W�7%q���z��w,G�T{+�2����񜛟׌�oB�zl��U��4P:�vV1��������Xʏ���wP�l0�\8�HU��^P���	 ����:)�։������4�y�*��gOA���F��_��p�Xr#��pI���<^����!��}YyGlŜ��fm���9ȸ�O��RXmc��� �{tH[eMGښ��z�
}� � �͈���Yu�XL�;��<�_��r�_\P�5����C��_*СBY���V��p'*y��iP�Vs ����m�����r�&����	�&z�2���Sw�j(n0P���C`.5�EnxK�X)F#������8% @A�ע�`������
�YQ���l�������&��s�u� �u
��ܓq���= 6�4�H&��\���}4)�p��Ҩ�l���~����U�z�ޔY�`R��m��+*'X�i�G	��8o4�{!G0ӈ�����7+X9lE�(�E�¸tJn���
�i�j��m��3���^�,$Q�l�w�6�R9�\�8�3z���(X�Ϫ�l�#��L��q���~`|Y)-��7�Oy \��[�=
�f�_.U�|�i8O�&Y���U��@+����
 �F���(pv�j�$�?��%�X1��x$HW�50��"Nns����,�~4�e,#<���oUvx�	��M�&������g��"�l��7�b�F�nGHj�]�h۳���}�9��2	a���w��f�S_�
�L�
o��K"�w�ɠ�m߲��pho�¸Ӭ�P}��DZ��g����a�[�a\G��RخL� )p�{�|�51������b����m��{�q�,%yݍ�jB3��u��U*�X-�9�(�hn�E�F\x��S4y"b�jZ����8N�w5�zA��k� 6�������ƪLm%�!� �� �~Զ�cy��9���"��d�m��Y�~F������0�~�L����9զ@����=��1}��cU��X�	7�T����d�M)���g{�(NB�e�d�n��6[`yj��A#��������g��]`6��֊�q��$�Y������(�ϛ�qoh�!�l���3a,jH��j	���
�a��a̩V�$.���Gu����~f�|F�. ���*��e2��ډ;%���w�sM���Ԑv:�C{�ju̶�A� ���N�"��Q�G7/��������T��K(R�YZ �TY�%�E]=I�w���R���֦��.�E��$��ut\lg%��<��G���Z��&A}ch.N�YR�S�x|�����/�Wzg�g��ْ�,�?! ����s堤p�tuN��>�����k�|�~�W|yGF'p��xJ�5���؜��;�n�X$A�����R�l�A��ſ�iH[R��o�L����?��X������fn���'���ۆ
�{&&��	��	�Ѭp��r����!`�����kPn(F�E��x�����>S��f�K��HQ��E;}K�d�w�2G�)z�y�S��?���C{�h�SV���S��nN�f�c�1��J�Fuk�[T֯E�A�XfĞ3�ZW%��f&��5�$�W��b����?�B�X��Y��KwO)MK��䦔'�F������~&�i���?Cu��}�I��};�?A��)Sہ���i�����pFƭ��avH��V/6�_���x̆���fYϠ���Q�GΙ*N+?W�W>�b��ڧpZ d��H�������]p�i�J���I�������td�qV�kK��cob�'�9��O6+7�6��%��.�~�����q&�rֿ����7L��̊H����@���
�mug�IN
<��2���~������qqF�����ׯ��6Y��W����z��P�-2-5��T���Y�4������L���L�Ɋ!݊ �ZR5�a�;��@K:O��K�%�������/��~S��ZS�����o	zsÃ@�}����!��#<��P�B�u�����U6K��3O�{��c�`*�6�,���O�Z�(5�Qwɭiʼ�,˖[lC:�
����b�]6a�9wʨ��C˹�QH:Òc�i�V�B�p!�f:{�6������;���$���K�w��8+̬���o2Xg���]
�S@)�Rm�!X̵!���x��o�%�S��b�lWt �6p�lX�{`�����d%dp�A.�)�l4-*�hB� ��LB