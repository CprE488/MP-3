XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k��)�Uƒ�>;��iD���I�0�q��^G�����N��� ];�S��c�{*s�?�D���`z���|�:ª��b���퐿����s������L��H���m����u��<��&/���cܑt�u���!X�*S�9�J�[+#�T0���XV�TM�Bm!s+�R�K�kF�6医��E� �ew�h߆�M�NP�B�I�|�or�b�ƒ�9�Ȥ�=����4~Fuv�͞�Ed�E��l�iYe�7hB2�_q���xz")�83�&�*:[-V�%�q�}[{@�EU�9�ݼKB��7D[�%y�}E�f;��b��)P ��=Q�i��.T�xX"��x�D$�Ǵ��.�%)$��6�u|��\B�(`�(FN��D^_��E�&���Q��|�	�᮰"��<`��)�z�tg!��I���4���O�����0�#��zs^1-Gr��q���IR��8L���#Tj9b��Sۘ�;��l��L@k70�Q������@rNCߘ�Fx���)KZ�g�J~}��4��J�4E6�.�B,.;��q�$g�Wȵ�n�d�z�M� ���|^=G��v�5�ku�ڥO�u1^�XD�M��D �w5��v������>�Y�,��KAϮ�ɮae���f$�R-ؘ�zRi�1�V�t�?���g�	Y'p� d6��jgr1�bOr�b6�R�I�
ųT� ��Go�R��z^�a��Ӻ��'��Q-�8��QiY�@%��*g�XlxVHYEB    1959     920k��9E#�4<�'�W�zfx�1��#�8Mg��B�+�h�v���G�Q����F��,dѭ��$]�D|Է�z�x�h�{��/�AZ4\=zJ&�W���`�s��xÑ.e��7g��Y�aN�d��C�Zk�,��6� u�+�0`V��s���Q�6-rDP��߶��Ok%���ʲ»g��i���8���4y2������ϧ��`N-w\�e��L�h;|��h�?��ʐ���Xڱ�y���0rN�r@2��͗.N�	lI�����T�2��j��
!|4�Q����1.Y�ٷ�KN�@��Ǟ}��f�v�ϣ|Bi7�K y�l�EË�Z��"A]r+�ݐl�$c�½��A ��"X�M�)��7�+��g�9���켇3��ӑ��A ��fŴf^#��['TI>NAR��ݾ�p��^����I�29�{���wE�{�߹�f�IB�/�y���o79�F?^X�sQ�]����G����@́6M踡�I�䏼U�[�V=�(.�(�eo�\>��q��Qt��g`3��ʍ?����Ҭ?��B>z���l�β�DC����� \mA�A�Ƣ��0Q���qBz�uc~����B��F��^t�~v�p��mK������۲C����-�A��r)��3����;)����դ���,�Z���C�<����q��&_f{@���3��q�h;/�BU/F�=.Cr�k��Ƅm��@�M����d`\��S�)�:��&ﻴ�I�Xv8�B� �To��B�^߹M�O'�}�J�f&�����.E�l��Ư�ҲV������ii���J1�"��n��CRk����F�0����Q����3��I�c��	�i�[�s.��&����*e�!f���p���٢rş�a���������m9ֺ�2��{;>�J��2_"��?�B�z���}?dٲ�@Ԁ9W�4>��<��
IB�\�Qq=FuA��3��=��a�ל�IT!s�k�k������s_�ܸ�A}��B���hPzE��mY�����P���@,l���N����������*�3Ǚ�l��s�=���u�^m3q�ͮoϒ}��i{�nIZf�J���[(�T��qy��^�#��]�}q{�t7������k9/�Ʃ_�l�C ��I?/
�ZV���Z�Հ]Q=��"@�VR���D��J���DG�e�%y��z����S����^��Tpr&�����\�mIU���!�2|p��8��[��2٩��/�S���� �]'�זȅՌj�٥`�h2��8�;!��2����#A	OȽ9���?!$��}!z++��ԱC-Y@oxi�3_#Yh�2U�m� '��	��&-פ��|daX1�͞*�p}S���c��J]�������o�U�\G�d��H?"�ia;bg������;=�D��vC�gJ0y�&��ò�}0<��$����
���t�z��g�,����'L�	b���p��}RWUKb�#�^�W�cz=nUS��$�	%N p�|��k�{ULFPt2�a�������^�(wo�8�����LjÖrV$o��2b/ei��K�<}Ц��y��b���\��AEP�O$ֈa�PoOٶ���$�n�a���d�!!k��sH��a���al�����$MV����q-�����'�O���ч������܊��g���G��/�U\��������؎i�	h�O����攲?�S��΅L��'����
�� -��}�<��ډ�H8��L������W!�Rk�f���Y���4Ta.˰�f,�M� }��Xɭ4B�����{��}��K�\;��ud�N���$���wjErܸ�ݵ��q�y��ߝ��f ѩ�L�8%�#����{��&�k�=�R�MD#g�5i�9r)�R�]ƿ�,�M��;L����k��U��c�����>L)�"��T�vǥ���\Z퀙 ��M1�ÿ�Р��V�kc���/G�v��ʄyMK�o�Y���$A�|�%z�WZ��Ƿ
�L�JI*⺛xu��^����l�jMwl����1�0 �
�8�ne�q܉��3�2��{Mܼ���m�K ����ʷ�i���{�i�B8�F��fq3f�&��D��fg�<��	k�x�jQ(��\�v��k�F�P���Y�V����}�9z�:�	t:Wf�:�������`�h�*��Jz�rb*�  9�d����S�f]��ң�ү��$�%/��>��[p�&I��sh���h�kej�}�H�tܐ��Yȵ�9�I��O���Po7�O�)Z.�f