XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���S"�����:_bS���s��r�XIM��)t�n�d��eA?���E�9��AV_��	%0�<-n!��H����v ��+7>D��}y!l0��^�<.�fz˙w�T�U@����&Ӯ�M�N=\]'�:�KlQ��sW���ɟg:.�a/t���S�ȏ%��?�/:��Ks�ߙ)�uvh�R�C0�U����2��&FrIw�&�Va#UV�E[e�>��$,1Q��x��h��r�VH���B�m)g��]W�ąyO��Y��U��Ŭ�DR'�
E�s��lA�;��\:��i
���Z�6�Sc���z���ۢ!0�Q|�K��_��/P�>fTh(X�J[��!�ϡ�)�MD�q,sb��X�,B׬C�GF���_bo׀���R�H���h���يg�,I����8z�����OM�T��p�3y �E��OGFU2�ZN�%�+�r59*�Bt����zoz����r���z���������n��Q/���Lq�T�ܟ��P�~�s�݌D	��t"�!}�� ҭ����2�q��i@�^���T��&Y��V�o���m�g}%�-���1����:F�%��B��l�2^����
���+�p���ۆQ�;+?�7p���L��W�*�I�	�K��Κ����xU����N����s#�x���e�V@U�` D�����}Z��L.R?�4r�w]�W�jJ�\NO�e'$�|��*vxF�O̺ЭX�gn`hp�Th�
9rB��2|XlxVHYEB    76a7    17c0�BkҲ�K�z/������82]�14����QA�����:B'�'�VI(�C��R	ߗH�jлFQ�c��@c��ߴL)f0�.��w�����'����3|��;�.+�L��O�M��O�N3!Փ��e����V/�k|����g��=fY<�]�!	�6P)�h� ��r�P v�8TQo%@Q�_����Ő��z�P4�/w�'�ȏ�2N�P*�:ʕ�a��+�p('l4Ӗ���O6c�M8�:xT���x��ۓk�5���w.4������4	T�i�ǌ�*a��va��l���m�5�Ez�# �}.���o��C�%k���I��Dp+D��aO}����/��;���\�	�h��S᮫_�4�j�E��K6i%����XÚl	�!�GrP��v�}<sd_���gS��P�%"�%[m]/�D��o&a?�4!���*�|5C|� ��pU��J��{�P��&5J��:��p,z`��a$��}|�˛M�TCQ%��p�g(=J�^���������*w�.�"�A�zn�_9�k�!������MTH%Ȍ-.��u���g8���[��� )x!�mNEH���b
�MMh\Co	b���GV��q�D��TS��+��~�_r��-n�y鲽ڼ�fx���W�}u)��M���4����Z@�܈�ln��$*������7��r�G��#�_�Z.�16����3쵅�{��,yo
A
�l�5��~���л�2js1o$.օ���.ѓ����;������J��y�Մ�=ߴC<I���{���N{�L���b
 .巑�6�a6��v�\>u �f��r���=�l~�]�Z$�}����!4�������Fz�0R`�&���a�2����������p���O�7'l�!��ȁ���*H��/��'?�����j���,]kcb/Q��ҫt��l�-!z��]�u�GV8[�~����|%r�k�ݧyK���yt-3X�e���9���Z�';Ĉ��z8���Y���V'�kV��?7���(b�()R8Ќ$�i�>�?_�Vy�����	9�u���K�Z��`�9z������{G&|%zy�*^�$�}W��XL� '�|�,���z>s��N�)�2[���!�4#��o6�lI�B6�����d�j�(G��`�͵��t�׼*0c:��y)�a���p�����I����C+���L�B	sj5�x��'���W�%�˻�D݅�ݹF�V�>Y<�)���>�kC⩈îg�n���U�,&�鄒��&*�Jk��{K�X����7҆�;競3"�K>�%��T�<��#%[��S;�u��BfJ�����P����0��y�1�nM\4��hy����개��&�ĨQ^�(N��ZҐ}a5ٞi�(���مK�p�J!�� �����Zb�Dмcm;<["�H����e�%�r���{,��/�鵔#՝������6��[� ��yo�H��e�1�y7�>>N�\pg}��2�����.�̳�~E�k���h6�L�����Wd7^ԗT��Y�o5QL�b�S��c�Ŝ�U��n���Nŏ";��[1������5#t��"�\D��kw���b{���m(xn�գ`S�zt�����F�N�o��SoB/���F������N�Y�����4p��r�pn�H�M�`d!%;n?tW��X40ca3�.^�
$��=9ZX�����;Y���^rB��RI��9�}�z�i(t�jc��	�O�@���\�a��K}'q�hۀ'�g���u�1��@J�YJ���ƾ��d��P�E#x���6ǢJ �b{>x�.Ok��_E��ъ�!Fʀ��%��"��l� j8�c7��-�*{�=l�|R�e]����$��\�m@U�  ��dX�dt<��L��0�*�-�b�FZ�m��VcL�x&8�����=�ݶ��G�=[~G����j _g�����_��"m\��Cp���V3	���#eH�뜁;��HX�=ֈ�Wn�B"j(�ߖ���7�]�o'z���0r����Y�Dfg)w�+�:��۱j����{&���UʖM�M��K��������^*�$]sE Ø�xx��ܘ�n��X�j�!:	�4V�]ϬJ�Ҩ�{[����3�I�{ %���!��fES��/u=�,8 E��oo�H�%��_j���d�C��%�ť� c	��E���W����-�c~9H���{6򖠦
/x��cn�A�vGh'f��}4{2����^�y)X����R�pw
�#��p$휞59�PJw����F�t���o!ʋS�\����P��ꌐ2���=4'���@��Q�;�C�\���?��э���e����j��8[�8���fhJǩ�E+b���;�F/ª��M��v�އK�����P�-��M��q�(4�J[��yd-���~�"���B��r�Po!�y�~��-E��3|���i�@�@��Z��m��51���<K3Ű$�J�NG0�%q���@��*�r�\~�A�y���$Y[���Qz/g�2��[�K�g�j��*�A���ړ ꑺ�&'�V=��%��G`m�xN)mb��%�'����լ!�A�DZ}}���2�,��ףW-�;�_dD@�N�!.K�l�� j�fU���6�N�n��@Uˠh`Z_�P=�N1��.��i���s���a#��6��uE�H�B�!�����-uѦy��Y]�����f�3e�ߙ+@�r�VN�Q��s��d3��D\%�P��ry�z(�;$9�*nX�  �*gJ����4?������1+��wP��A������׀y$�HV,'n��M��I�2���� #��I"J^.��0�OVV� ��m�	�<���p>��4|Ұ������+�h�1g��HА0��G�`�?��:6���٢w_*�^�B�r��4W�P���s���%���"��u�h������ m���b̲���K�=b��yT�O�pϔ�ߢ���<�(Z�4�$_&���ܷ*\��z4oˤ=���p$��p��+]��CK�FV��$��	���M�Rt1H��v,�`�<�U��k��a�Z�m�ͯo9�$iOT����v�0ec6&�vU����I���7X�`\���*��sV�H�RW게Clh��:�D?>1c���'а�K�$�/�_6�.1V�x��[6QB��5��Y�n��g�����#����VzLUFk3m�q7"�ʫ�b��?|Kק��b�U���P��9�݉s�JJr<���j�+f��1�������\����
Ϭ�A��wg��ũ8(2@&q�Z���婉y!�˃�be �vJ�����[���VRǓmob�����*���y�"�MC���˪`0F0�ƕ*s�vV�^��0����¥�B:�4��I�1dp��!ͼ`ggWk5�)Q�5d͛���ͷ("�u�X]0υ��2��U�w�y������$� �%��:�g���mχjݫ/$,����%���v�e�z0܉<��z�,�+�wNl��!u������^��
�8�W j�³��nrI-n��MqP���7����+r�'ŇE�Y���5ˢ�<�=���>M�yH��Q4>��>��e��dz�ȷ1-��L����z֝�#��G]nWQA��=�T	�
�#�'I���p�%Y\q�hݤH���=��H-�V����'e$��7J�g(�{���>�;)dy�L8$�g���%X�l��8;���zd��+�2D��t�?[L S��,  �P��+L���X8��l��cB�Wf~��{rsڸ��.Д? ��guځ8���iXR#�?V���P��8���k�|�-���8Ԙ��}�i[�����z��u��QW���FWi0ֹ� �laF��u��0M�������8�_��s�jط{���Ŕ�hF1���}G���2�H��Q��5g�R��^?T��Ҁ� ���Z��\�N/�᤭|%x�z5�!����"����j��oE���c��C��
�	m�S0�����Z�5����/aw��<�e���_�h��7����#?�6I{Q��?�QD����Ar���/ӣ|�Mx�@�sQ�R{�L�M��P-���bi�7�W�~CTI���r�j�(����Vxp4�ImʼV���9��ƅ-�m,J�#-'�J��).Pz �ݪ�/�(.��P�w�ɟ휱�4U P���_�e�������J��Q�:���A��J��^��R�/%)��i�G�D8�CϦ�D{�[��5\�eї�]�:�]�)!$�wJu�7v�ƌ�����pN��{y�fܛ9��3����YmNK�h�q�p����v���������bp�^ ���LH����L=wC5�������w�-=�_A����lfN�`�Ɉj��Om�o�~{�9?�KT�=E��� �uJj���0�+̆G�k����QY��Ƴ��x*,
����l�r��9���UͿԥ_m*�NZ����x��n��j� <��COF^0z�AR������E)#I�ֲ��Ю��4?�2ӿq�O���S��߄Yf�饅|!�����Ь�B��,���֡r��|�Mypb��#���r@Q�z''�j�̩ց�5h/�Q
:¶���EA�C*"6)�x�7����E��E����
�	?��I\�A���r��E8\�Ҹ��x�� �u�oq���H<�?;��J���ڕ��Ɋ�-b�S�:�z��K�����J?"O#o�l�|m���la%m�����:��G�x�*�	y��:/�B����"c6��X���o�
y����4A��\S����5��mↄ�/Y�\[���2� ;&d� ����	�L�y��`�)����Q ��ٺtd�-��Z��Ӄ�8j�p���k��]qh�H���a 'h_o�M+�
�.�Tݜ���l�.����{$_��c�N���<�;K���#�KT�ڨ>�}� S��<��^>2��M�WV8!�@�X����SR��M��x�m'�Ƶ�=�N�P��CsU�mo�b���P��P�i�b_Ϧk�q�܍)�}�oS,�<TJ�XL�a�Ӻ�3H���t��O��مws�zGDC��|	q���qM���)CH���!)LtU�ciU������r��0������L@��ݕ�A��H�q��1��wvomGI�Vg<�N|rZE�ad���j������䕆�Ķ��$����۟Z��&��c�6C����J8�]���D��T��W��}b�C��p � P���b>��{� �^�`]?_ۣݔ�a��Q��.��N$��r�؃�������&L_�9�p�TI��Z���bJ
����0F��F<=�����=����8S9.�z��S��=�����hHH����ơ��I�����߶�[�?0!��l��QP���HJF}�&{d��u���Nq��t9|�Q����Y��<��å��
R���'5f��Ԇ�TԂ����WFg������[*'�����"a ١���m��C�j���e���}�Z��;Z??���b����
O͞��p�L�wl�oԗ���-���Zk�m'o�S�`�
�6�?N0å�	�2�(~f2v�U��RpѷA��%�-	��x,�ˠ�\8�g��C��2M�my03�4�<@o��t��R=}}�X58?��p.1����ӵܱg�V��w��)�����,���i#5ܰ+�m���~:�f�o��i��R�f�lo������A�`J��gW)�!e���<�����D�b��g��5��1��4^�� ��=mf0$:(��	+{y��;h0\<��g�5O�RֵL�yH���Y�� }�P�p��)W�*�  wtO�1� �g��{Pȋ�w�n�|�{�B�GbϾk�W��#Y ��;����