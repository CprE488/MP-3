XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W�����K"d����A<jP�jK�S�W
;0�sP�q_ �`�FrW����a�������Јy�)���pMb	����3�3�e�iB�͈�&u�(kR�4�]hV��k�eA��W�F��:PT�����5�-SE��;���_H�뱟tl�����X�+m�}�^�����j�V�Ì�ս��Ш����\+d���a�c7�3�D�?�?��1/�zQd:�,rd��<IGA���� �k_)u�:�Ϗ��2ƥ�/�,]=�u}��j1mm˨��[r�-YA�:�:R�.�g�r���K�n��?s?�	�e�{��m.�;�A�P
��k��ʓ!B�1�%!zP(� �2��Ō�W/$��`���ˉ�;"��Ƶұ����6IK�D�H�árY�vL?������"����������ٛ����@�c�Ѿ�:�r�<�@$��%�u)�:�q�iƈ�J���C/�P�s�e���� 	�r��2%�������|M*?V�$���B�#|`5�(A}ڢbċ>���3�-+m�x�c��֯�S�3� L�W^��[�^w�pa�yI�[l����J��kNßF蛲2�`�����X�:�;lR�����,[��FP�f,t�M���v|)��8�V�+PK�$#b�,�<ƈ�����h��q�4�} �A%�>�����g����7D��hń�s���f(D�"Ft(/'+���Q�*V'�R0��&���&
�5 s�z��/pX�X���
^��XlxVHYEB    3d43    1030�E�&���y�YGFx���!��p��0�M���)��}vQ}���Q��;��*@�WǷF��B�wٔ"z���6e����Q�/N����&��� P^I
��P�'Uڵ��ē ִ��#�t�+�	�K��~)T���'�6�#�����XS��CY��YBmzAʢ��.�ؠ���t��ig��4Ŭ�1���q�>W6F~�cpo�D�����R�М��@�ӌ�`�l�wi���&~,
D]�6_��s�Q�K�CO늳X񈸤!]����)�&R.�Fh�v�P���7l�$Ծܯ:/����������IR6�O�'o��b]�g�7��/���S��ٿ>�d/�*^�H��I1rNu7s~iW�
�u��g~�T�uW�{Y�k�Dv�) ���Q\���8%�^K�����)Yҏؠo�!.�)��[R�J%Π�9N�ß{�l|ȆV�4�m��E�,���@���2k�r�x�@U�m�X%�q�7����S���^����c���r��y�<��/�ژ�M�%�H��1`��3c/"�i���C����.~�ܤW��#�YB��ME�}�RB�����zS���l���~8���Иq�E�j�_�!�X��C�x�1�k�@�;d.����J|�� b��µ�R3���ROo�ؤ.���ęMdt�a��k�Vx����<(/�]��E��O�:кd���*R�&�Rj�V�����3��Ƴ0�l[��Ifc�.i���E����N�XZ�ޫql$�iG
�e'ձ�S�;�qB�-F8��TS�Q�A���c�k�����)E�c1��'��SӇ��2~�	;���y/L��O��)��k��G��皦���U p��St(��z��ՋR�B�p��㣉,y{�-E��^��[�*�vB��e+���	
v��;�/�*��cf'�D���msF��D9)������/����֟��z�}��q��|�iS����8M :|��[i���K�6�]��ş �w�B���a��H.���}TT�.���)�j�z+y���z���K�Ӫ���m�F�+���L^��ߪ�V�Mj%�XzG���v}f'����|��-u]�4���0S��E����6(R����g��W��3�e���0�����M��^���@�,���m|��*$!G�fL*�Q?b�|?W��h�U�E?5D��;������ս����! ƚ��iֲ��yy�رzeo­S܈����\�����r�|;�HbM�b���V�����}��Mb	�
�R�
���#;��2Ky-��F���$B`��6�P���t��K%�G��l!4࢞�>��ŧ���D����=�Z�Fa-��Źy8�&�a=���_m!V��KW�����T�~���)�87m��5�i&�E��2��[YԄL����O:'��&f���A(��@Eg�O����3���m���s�_�ҟ�������o^�/.a�{��}�+��]n|�t�O�����*>�)����%�R{Yݔ����z�Y��V���!���!�,�~U����q5�<KZ�p�{�Ag��v��w�q擠7ۛ�a�uB��o%�mll�xڊ�����w���
XԀ@K.2Y��������D�R+�[��ujQ��~ ^7��
z��1���S��n����дe�W7�6J� F:��3g�IX���4<�.߂*
�<����%�MX���l����k��{�n.����$��������o�������
\C:������������욬oK�!&��D���"��Gd��,�'jK��VR�
��aeP�h�7}�
�Ї-%Չ9̶&]��w��Of��E�,�4q�B���/��<(�e�5�"'��FP��3lf�Y�#F?	B��T0:�7��   ��uE%[�%��1��)�;�>�U(�:���@K�f�_�.�wky� W��h%�.*."�@�([	�9�%�h��aP9���;�0���Q�5�X�r��VvR$���v��{�����9�ȍ/f;c+`�Q��Ч*�a������c���gC,	��u�"�:p�=��\�\`��A��J(A"��Sى1t���ʵ�F'���c��c��-=�C��.6�x��	Dd�!��.�Ep�k;H�,�M�iϒT�����,��e��$�	�a��.s�j�����P
�շ�Y���ރG�9 �E7H�5iv�Z?a�C��������/v+X�*p�=֍��N㔣'տ�iB��Qy�!<yYx@<�,/K�2�!T�X���S�w9qw��i,���Z��_;X���e� �QDҴ^t�_��L�'�+Ğ�F������.E�$�B�l!�M���W,��3ڶv�K�����Kp/1�|=�8^����9ʍ����J��~��cҥ�ksW����90�i����޹�X��i�-{LѕI��L�|W����_��`�^qc6ր�BH5�QZ5H�c��W6�e�[��_Y��8x�����TJ|�a��:�B)�`�j"Z���a���C}�ݨx�9D���(,B���
��Aݟgp\?ڷ\��������ު� �/��ʟ��L���:8��']��dNX���3�{3�x A`,Q�i���J���B]h�]t�6)N�-[$J��,�=)T�j"P�1��O����Ro�8��Y_߂���C�uU�^u�E��<��iB'|���*��!�͈׃�L�bR��u�H$�< 5D�sJ��`�w�8 .�/E���zl����7�9P����!�^R�{6P�V�`���y�S��6#{�ϳ���6y��N'=��}�L�|z_>��O�,�A�/����R)��/�)w7�OZvT�e���z�P�<�ĨV����I�8�%p�\�1�� P�&�z�ע ������l�&rZB�'�D���p����P�L.#���aN�~�!��
p�_W2�ts<�u�Y��[Q���^�����mbS�vn�%SY�B�p�B��zL��QLN)�>�i�"Er�a�H��(uY��g�q���N
��w���hp���x6�r��tRap`�d��/�^�)�'���r���g24/�0{�����8:V��5_����P 鞏��Bn�A:�E���Rخ���������n�Ņ^]��[��7�@�û���^�.�ʬa.��?|r~� ����Y.V�����FoL����w�{y)d�^;����"!�����8�U��Ԃ3�&���NH�ˡ�ђ(�S	�����o�?~hÆzQeQo���k�'P�lSe~��k��B�<���� 5u������*�O�YB>��{��C/Q�D(pƫZ��[����5U��>��q7��2/����]��u�)-~��aa�'����'�����ze��N��oՐ�@�9{i^T[�F�.�����yb%��q�� �>�X��:��#
EF7�s��r(�^7P�����y���3�clu�Գ�!�6��G��9:����9% �)���<�W�-�:�,G�"G
L��W��ޘ�G@����0T��n�����=�� ���� sȦSX����^7 ,�uݨ�Ɨm�E}�QVA�
(k�*mNЈ�=����̤9m�n�`�_�E�-��"~�q>��K�-0��������6�.��"lK����,[4%h�*ǎ�	�I�;n�\��U=�l>��������ח��Gz���@�O»Z��i����q�G��@���
)A<�0�=뎸Wd'oJ.�$�1P�ۢ�!ٖ�	���W�oewOtD�n���e�ZEᝪ�le�/��-r#�6��y�M�	 i��NsF�iШ����ؤ���;��uu�/�E^e�'�-�K��&���^��Uy�E�C ��p��R�AO�Ь 45�?ߛ���<���f�nƅBnX���^8�@Ň@�>���6�E#
��w esBGC gR�D8P�4�1�C�����(��ì�cW��M��\���er�z����i{)sЀ��n��