XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��e��ÒI��.f��H�_̆`�U��f�r�&sЮ��g*
��jp��t�	L[�܈���e8ȥ��C�Z��	��F����P�̭����$�A��E�@���S_Y2�R[p�Y"�G]J���ߵE�r`�Z3����᯻��$tꎉ�EEc#�9>�&����&��'{Uf�*�3O
�2L,���DZr�=b.��B5�6sLq�a�����+�BL�q\�Xj2E���q*�2�����՞�m����q���{\�QP�e�`��D��A�>-�-��G���$���M.$���ZQB��q,T�?E�\�(:E�JۉWR�HU	yv�&��d,��3ʭ��z在"M����:�k@����U��k"����}�#L�T��I%��uHϘO�9���RѶ[P~�W��x��c��yj�<cckJ�~�9�"��*ۺ��4l�n�UF����c{�-I��y&u�I�"�5�G�ͨ�?���r4��:rܳo�'��6��A]4�S􁚨�U�W��M==�%Н�P3������į�"^�`�itfu�cH>�>|,{٫_Ν8"ԥ���l��mⓒ�}�wZ�m� I�i���VQ�?��П���[�N}~��%Y���d�d�4� r�у�|*�_(�`%����&x";*�0�������lq����l��4����-S��tW�T�]�1UwgK�䬤��y�!ia#�b���N�C�� X\ ��f�������钣x?:�K����)�o8��ތ��XlxVHYEB    1959     920����>��dz�l��1��W
�$e<rZ� }��?�̏v8i�������bE��E�G����_?�mg�m¶���b�&�sc]^���݌��$��Rq�4���r�O>8�I]5�l䤵��X�
`37�|���H$�e�ȯ.���*�^ႆ�ͻb���K}�G�.���79�"Q���),U�v�X�QO�7���}u�.��xJ!B-��x�K�|��D��@�rEKnP1�#�/)���N�`M8|n���;Oλ�9�"/��1k��R��6|��5�ڶ����: �6�A����Mp<}��0OP٪��\���*�ӥB?�Lgç�'���m�)T oE��JĥE޵�����%P��z$�ư�!��� /F���l`��a�·��5���O4<�f%>��2e9E��,|�yU�d�TϹj�`��|8�M��x���R���f~3 ^����#�r8�v��0��uO��s�I������E���(�܍�.ٙZ��;��<1��P��;�3�ζM6ӂA�8y��02R�>���4���)��޶?�6���_� +�{!��	'o2k���p=AWd$��)��݌��H�^�v��5Ҹ�2Y���R�c��&�O��;���>��w�cb«���mS�_�[{<qN�����{~r)�-���tD2��]�*M7�&����dv�m�5�f��뽂�v�L���>e�����\R����	km������	��ǢIvB)�����w5���{5�8�xq���l�3�|��eQ���Q�>���rjoA#S���Uv�*Z3�cK�	.�'2�p�[~�@�լ�2���nK��ۿ<�3+]�0��Bܘ���w�Σ��`�����97�MH�Uw���lC^�����8-DA4�y�0����]��9U�`�#]k�'�W0o�@!��eK��s-���/
}'>8K��av[.�m5��aCVZ�V�\���ט��:����aծ�S
�WK^e(x�͉���)(7� �C�i�(�󩰊
�9P�$a�5� w�2,mOK��z&v�!f�<ɋ����<X��&���<��1�+F�x�rR��锿C����b�yS�jjs@�V����Ist:cа]��Z��Q���h���q��e?}�9�ŵ���(�@�f���G����k�Q
1K�Q�=��Ǧ�!4�o�m��W,sL����{�"�ܑ4��\I�)/XoP[$���O16Rb�>U���ԛ���Fw���[Y/<t���ȓ5Ɩ����H/S��xpSG�Ȟ<m{c� �[T�䶗�}C"���>��=a�d��!��=h�SG�!/ ���7�"�\8B��]}O�o��O���F��? ��@}�~�H��փ��j�ԏ����\7����� ,EA�:^}m���*�{�{�������b�@d�O��㻃��@�T�zS��-6=h/u*�9Sa��6�)�{���@���̥|\��Y���M�;�G	F���2x�������g)_���*!��j���cd͜�
�Ep:`��0�Ό��U�S��ްN��Y�K.|��<2RG��]w�A˟�)L���	i96t(�J���9� v�l��2�~�WD� t�	�z��=6�2P ��Ϻ��,\�[ì�����;�oE�Q
XL������c�f�</��;��xu�U��@�a2�[�~���'�B�՞���B�k�-��� �k�1�<)�rE�'��)- ze��d���5Hc�ꧮB��pR틖U�����d?�k>�\�+�쏶���i��c�s}�L80%'�:T8�s���������Y�:��0?�'�q1���qs]�qvB��J�dF�7�y_ _�\;Y��&��`,�u|��v՝@s�E��̞ ��Sn �)�3�0n;�{f���z�;�/�g��\1�C����bW�N�O��׍��$4dH��Q��p���[�|����N���+>���t�K΁���o��x��R����O8A�E�c���b�Ċ`�ܐ�65S0���-.�U�W\UZ���+�-��Q�=ag>ebN�V)"�_AtMi*L��6·����~ T�y��_�S�o�j~o���=�:���T�$H	�roU��L���������Yv�[k����gG	L�Į�⭸��;�H>��'NP��8������ʑ2��fT/	7�Aˋ���[��n^�r/���,�4f�d�(R�Q<�K�f�w���.��#-
˪/�ոsJPtb�I�g�1\gYŐ�I�q!l�S|gg��<�t