XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����/�5σ��f�6� �{��p�\��~�#�=˽j�a�fx����C�:�򔿓�kaꒂ�6\���y>�Jk�}5����ٔ"�&X�Ә�/�`΋����f�7�d]�d�E��*�6���EԒ�GVv�{*;�m�<&�bܠ%#ph� ����ȣ !�fi�n��](s"���K��.r��w�Τ�E��ξ��;L�"up��7��Em��~�i�I�io�Y��#`����{|�x���9���5�������1�<���i�^
�w������sS�m��Ɨ�3�I �&O����甾��ZEv3���TCٱ݊}3��g��BL�0�]:o�1�KX]_/jQ�[E"t �c��]i�7<еÓ�t��A�O�l����k�k�Pr��B�q�Oט���N9r�b�L����_����O��62���3VF��9I��U��qty>��G��\h�$`%|p���%��k�W6�5G�$ΈuN���/�e��j.�%pL4��F�+-�Bu<�xrf�Z�;E�R����Xl��FL��0R:в&�a��_ض���n�kH!M4�_� \׏����&����o�&�ƭ����D'���#�:ȿ�|�����$+��|V��g���8��5�@��R�;�]�-FmdE�S8�Y�]�4:���y�����h�����z�S�W%�,����N���9��������7>{0pS����RM���ʌs�Aq�G}�{�*�F-����`=�XlxVHYEB    5e2b    1530ͳ*���B9U�[B~��G}ѧ�
m9�%�X�cx�}��X�	,��ⓖ�%wh�p��C��出>�99)���N�k�|?��ّ��u�����Y9:�H��մ���GVf�S�+����e0�_�'9�<�!׭��J��G���� �7���Ej�%�׊y/�ݺ�a-��\1"�$q����B��°0�A��F/��ң˺�+ڢi5��NC�������:����/�y��8y�����L��(u�Y���zKF�" �.���QI2^���髐��A�q�T�,p����Nη��I��e�'ː�|�ĎF�R�u�fٔn����;�O���πd�鄢���ZIS�۔��ǣ�:�r�V�o__��q_�/M2����5��`�:Z��ZS_�����
+���Đ�<)9��t^�E7왅q'#ާ��3\���<�ABLZn:[���oQ�7�M�Mr�9��PE&أ�
;��ǣB�W�V��ã�>û��܍��=RVH!k�X �HN�u�� ��i0E3����*�X��V��\��i���h!窹W�)��r�`�vl۝��.�ЗT�1�\r�d+[A���+�H0�,�g��rF�ɴt� U��k�~w�(!A"�X,%���&���C(] �)B��d��$��������S��ڋ�Y�����+��랆Y��>��fϼ���4N�������)*z��F�Z^�"�qy��+�����W��>����<�"���ߎN_-)�����,Ш$��%����T���e^4�ǳBD�҈@��O�%����mT����P��D���j
<���"	Nݮ3�J�=&�K���ƒ�e�t�4�hZ�S��������������|�Ϭ�A.'RI�� UYR�TᲰ������+�R��7e��k�jVA����-���pK�&.��<�C[�= �[�F8�i�Ysq ����7��f��G�_A��-5��<:�<�=8���p��!��e��梾�n2R�#J��dȷ�䁐*1���Gv�ۺ������2xZ�J���,��GDӺ�m�� ��9�6�S˘<0BSq@���8�^h3I�.};JXs��
�����(L쭧=|t���?&R&%i�H�l)�*������J�f���G�c�ϴ���|��E����EE���^�qA&��}�M0k��X|��ʄp �Q����Q��P��k$�Q�h��?�&l�з,�����ku����Z�l��[Q|Q6�R?��q�z7f?�m�sTc�9��﹌��v�ң�(���ϋh�g��Ƅڏ4�N��A���Y��v��V�Ox:�28�'GL��^�9��6�"b���D�)Bf�nK'Gϱ,��B.���N���Ź�Z��_�|��h��^s]i��e�Q�@���>�'�!�h�C(�I�h?���#��>}Ƶ��n���(��`KT��J���ջt���E����֊�XB��k��E|:\!=�g�Ԙ=Ԯ�`Ä_"h���]�"!S��tE�2gD`��L��}���X��_��-l��e�[���Y䐪�N���O��.a���ڡ���x����� �㈷z�x�}X׏�2�N��>W��\<I
�X�v�P������k�&�� �����㨒#B�[���8}/dL��8")	�Y�1lP���ؙX�ozsۯ�P,���Q'�	�vD{ v} �4�UԄB�'�P��������_!�0͔�E��=͸A��8�5Fc�h�_,ǪQ7l��B����lU[)�_[�)��?a����Q��#�X��b�0y�r��"��}�̑R�I7�8]�
Z���c���}�wL@3�������#]��?yeOb	sT��5�(�9\S����ꮡ<V��D��D�؜�8;�����E��W0}�������/~�����kV펃���pn�c+�>��uCDо�sSn��N.�$x�O���xzI8��g�}g�d�Bڡ�%ipM���1�;��z������Ȱ67-�d��$I�vS�r&�jrl���i�DG�h �X�6�Mˌ��.q=(8��Ls5�_��&��>h)��)�^'߱)v�y��*F�Jt����$�kM���8��<uq8�U�m����r�<��w2���`T1x�n�NӥuxT�ޗ �_�c?�� s�E�,4��]���{�ْ��`�tzm,��5����~�W��u�U�x �S������`8���Rh�(��E,?�}���P�{bW(\9f���	��j������|�^q�|�����У��}
���;��g�E���s@C/㈾��j{�p�AMqbH�,�t׸�,e�X"�1)�EW�L����ձ�5l��6�j�v���P��gn���+ n�I!JI�}óX<�7���sq�*�~��U�M�`�Ɯ)�$07}Wܸo�1��X�^�F�#�*��V�u�&��H�uiV��;��Aj-B��Nhl'V�!��1�%���v�:q��� UA>�;wy���F��)�D�o�2�6��\a��[>��Lx�����B�?���db���}����W�m|��P���R~t�m!|���Oڰ��"�Q7�@���F����N��}ҡ����v�A9��3�ai��gL�G�M'�R�~�v�y�R�;�uGH|��sް��K��&T �Ք���ڶ8Li�W�������5�dۣ�	�1V���/���5Y73"�SS@|V o�/��2�"T��^D4o��(2x�w��遻`�'�������0��tRX'5�n9t�c��Z*&ɲR7�K_��M�Elս��]1�矃\���`T��������\��§����,A@�z��-3��*	P{j"��}2��3��Ω�~�w�H@p�Q#}Ŧmt���W�����&�أ�Y
I�"�̯�;k1��.v3�>e��˃�7��lY�����C��D���һ����' �&q��"B��T�3�x��Of�x6�@(�����6j���6_�^��O_��+J|?�qF`92���*�Y�8�R 70'"�H��o��k4�Л���|���ajT����}�gҕxO�W�dk��/��FY��`�����=�i��Y����?P �  �i	�m-�o�w}EVs��1C�#杣n�
f�QN�O#v�_- �zG�S�r��z������L`�;Sf>z_���Oڼropz��urM�.��4m��u�/RJ(��G`�5;-:�G��g�m�(�g�mq\�oq��g*-��	�d]�%�<$����Q����'q�QY�	�V8����P�tm:�S�rbf�d�5�W�����ٯ��%Y�soҘ<v�}���������8���Y���'�k0��	�~��B�7���⪖]�ˀP���D\�� ~Ks��*�q|�o��`�mׇ�s}�]���ne{�F��S��&�d�Ï3^���dy�c����#�K�l�AZw�&k(��/��xS�*:'%�ɦ�=xj��i�g��)4WzJ��+Xu����������x�G`͍��.,����By�T�IK,�͠ȸ��J����E���l�q�}̀;}*�c�.��C1���������X�"�"1}Yߘ�~��������dz!���P�P`͗�]zj�@�o^�L��S󲙬�z^d�[�
��d	ַ��j��:��}�>�c�ݥ�Vh7jcz�Q�)Eb�<GR�C�ׄ!h�|Y��2w�׳[���vy� ~b"��Y��}�߉s��нp��x=���{�A��������@��aEW�7i�Z+%������!��5��!/�Qi�au�#�F�RU{[�u�XFB�����7k+-�����}�F�[kӛ�+�j���M'xm��#���yi#�0�T+�ZF��Z�x��s�g7���5X�Q�Jٸ�o�NL����NS��(�z�S��ǘX�<)�n� 5���tޝ�
��W|�r}<�\�_�%�Ė�Y����m��dh���Y�CJ�@��M�-z��+c�P�����e7�Q-Y�崻�o�4��ihG��0�+���T��}�F:�T�vn=v��`�("dѩՓֻ<b�ˀ�1�D;2)��{a����/�Pw�ovP븚h�7ֆyJ�T������i]�?�g}d��s�lr�3#UY(+tqƽ�bR�!2&==���
�����h��7�?̷	Cُ��W�K�MC�g��C�O�iyV0��%$�Mjzi��Y˴~�2�&&w�%-��H�t�@�E��]&LԆȱ�I��r!���ሉ��;�C:#eb,�\�J@����[Q��������t�����aj þ�MV�<�6^Cm�h@Q��n�|9�������z+m��I�q�S@�םn�/u2b��/ �o��GB�TI����ak/�3��u
�sN�bP	ڕŏ�s�"�fj�0	=}��MR�2�e8�-�t��a�[�'��������־�D�B����<t�w
�l{��z��͉�la~cz��g^n�^�����*�D���_qzz����v�c&0_�z33�]<obh�oD� ")���i�@J�O�W�-�	��qr�{3@Ԇ��,�LB�j�qn neI�Gk���r�ȝ�v<��W�hD�\U�-R|����c���_sѶL����*Lq'�7ҵ2�,�1�}�.��c��{���⣧�m0��h(�[���)ˠ����3F�z3<د�q�D����#cQ�Օ��B���l�D���éŮ.�a�C�PHx�G'���=!���#���8��YUlc�$����u�u����י��氤��r\���D=�ܚ����fP��帛#,i�I��o��6dW��%9�a�ܗ��}���K_����FP��q�	7!�jƏ�P	���71'�����o�$ɧ7rW�D|Z��ۈ�Be �Q�}%��++b�g4y�;�8�ܞ�����ē�%X�m�8���c�S����J�'C�~�m�&[�t�CM`��;h9����Ez��/����P�p:��R����³	>2��P�����r�ٷ^��v�:�9U.k�!�=��ج#E��D�&�gQ�~!�ǧ4�&�� �e	X�QK}r�����Қ�Vں�T1*�J��ya=��}���v�}ĸ�����(JV/~d?9���������3�wN�ꍵ
cTuz/�,�F��2P?��6����dS��k]���I�x#�c{��j��{=�(e	��kgp�B[�9��u�y���N��/0�T F=�N��J����9`��r�lE�q���<"��j�hr�}��ϵ