XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���{�+UQ���L�kв5�w�Vq J�۽�A�eƁ�I�dt����mM��r鷕�� wR����jK@G���zӬ���֘̙�a�q�Z���7N�}�yrnB�K���5k���죺*�E�MA��cH����_*�5�sa���WQ�k���#9�Pp��"���c���Z~]ୟ7�K[�{?�'�łe}Б��*�z*S����}�c�t�R@�����!�4�8�Bd�9O<8�!�<��e�)��H�����JW�=����Dkf��W. 
Ψ�u.�sR���,6�4���}�	������^-��+cB,Җ�j���~�b�s���j+`�ӕ|���2T
����	i�Ш߼y�y�������H������Į9,u�R���f4{%F��
%^A�L��GϿa�mw��K��f8L��F��wφ�� mp�.Q�������P}�y�"L����)ǖ2w_�c�w�JD�kB�-2:۰��5wz%���{�����o�c�hh?Z�Y�ۃ�i���gu�r`~�<���\�wy.M�]�bz�.��MyS�1�I/��Dw�d�茅�	T�`-Xp�j,>�CʻJ�M���d�5���ɱ)q����毨��������� �`M������?\�aV��~p� �l�?��6%�o&6x뷭]5��_i��s�'>��b-�3I�rx쟽7��"l���^�l���סm�@����vkQݗ>XƧϣ	XlxVHYEB    1a2e     8b0�l�f}�>����e'�]\?�#Cl��pX!��i�'���B�1�,�"�%�o�xU����@���ޗv�c��V�,H�vOL�w�6�>'��1�z� ��ϩ�������@Ԧ�cA�ðĮ�U��q0�S�����������;�%M���~E�h�7:x4T Ŵ���d���Oi�5��g�,L���&����|��9�Q�/#!aa���˻��������>@�6e'J��ֈ-�OƲ��G��~��&�x:6krX�eΠM����jC�e���}��� ���8d:���M5?��@7���"�w]�Y����9#k
2�B�S��#e����76�9��!�MM-g�+1qV2��\&��?I[�{&��A�1�w��J	[Z�S�${2W�iy�2�d~Q�fO��Wt'�sa�'��U���h��E7�P5�� ��H�����Z�H�D��O��C����~�Q�4��ه�hr��(�I򆛞]�2t��ϯV�5���S_UiqkȎ�<e�*B��!φS��T���>��u��d��R8�~:��8'�܀f�lx�A�0��πص����T���'�ڢl�R4���MT� ��o�/`v�X�Ԛ��ŀ6�A-;i�_��\D#E��C��8`�m�i��E�z*��Y�M�n��
l��l�0v6�h{F��xĉ�i�|�y��ߣ贕������������TkV�q-��c�D��Ct��(���o��Lc�	�^�A����~�0�ױ�y�����3K��lC��Y5�B��u���J;�0�rh�n�Őc鵏�/�=�-�x!u^�e��_d&Pr�H�.O� FhqfX�$���.-�z�}%�9�l�����胯G�F��4q����ą���܆iw�V��A++���A�Z�d�#l4�|�8��_!�i�վ_���_�9�H <�Q���p�9��w�H�o���'n��c������Z&�9����3�u>?�3�h�}���)F͙{'��Yx�ʼ��*A�F`(E>Ư������zI�i|���]Û����]0t�a:f(��	���^��7"�mdE�rс���'t=�!�q���i�V.`���.�u�HE�ƹ�~��geϢ�����i�����{�ꞦR��K���gcv�����a6��U\k̏ �vM0q�MK�ʗ��-V��K���v;X}��L���mc�s�44�e�8���p�7��Q�7\��a����}�D$�Q1*x(�𐼮��mg��s*�h����,��o�$��es.!'�z��+-�j�S�/���w������ï�Y�N�0��� ��H��Q�W�3m�_�r{^����Q8�h���!��� �����B��2�x��kM)�%`Tn��M�o'�}��agS-�F��{����0������	�_����wE,��:�o�}`�C�y���Af��@˳j�hgE0��Lth��!��,�*���B�Y�D�����,���w ���$�h��Y�{�
~l҅�b�/g�SF��^pj��N��}K��Z~��e���\�"x�Q=8���G5pz�bp���#�SAz�� ��W|N����Gu��N?KM��6﯐��r99ΰ{5�K\�{�7��^v
]!%�Ol�Wsj�_�'8��@CT/��$���X�.bu�[^|C�I���*a/��j����j%a�mA���>�/��΀������v�g�CI2[yN������6��c�>i9����c*Ea��T����|�� \��2
�)���bs~�\�m�#f��SVA��ʈ[9[J'9g4��l�0�D����~5ޘT"��w]}���F��_������^<�k�(�$�0�hō��?�����L��'?��y7��<�J%B�Y�i/��@Hvs�#� �2Ŵ<��T0g�3�3f���'�=6�ۼs��8>;��CE�
�@r`�z����,�<�>N*\��l׶#/���芳~Թ��<c,�7�p�q��������������/��C�Ujx_��i�w��Nt(�FhYS�\��9�,��"���nC	�T@�vH~j��Z�
.�w�u%�e��&��j��S��A�T�_`���%��[̤O]�4\�D��B����X�Q��<�$������z�F}��:�A�%�R��L�@������97^��q