XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^�ޗ6�*��cy
}���S1����~��y7�K�-?&���e D5Z6�N3##����?N/�]�'��7y��Yk��$j��bi����V|�M[a,ݒ�D�o����W ,��M���a���Ɯʃ�>st$v����9J�+�r�G>�&LkV*�-]�L�&���y��2^/h4�1l+�ʰА�Cb޲ˠ+���b���$f[1w�Z��j�M��k1��ȫhl3�V/�E��U!h��n��2\�;����8dm��W��kD?q7��#�7�	z�E����a����ŧE鈓��G釗��ǧ��k�k%���u�>h�)����C� D������[�u�&B|��bjD��×��|��d}�F�n{#p���+�'�^�2fƕ� �>γ0z3Z���d�uq')o�M�Ml|���֒n@D�Ϝ*y�-�}�4]>X�dȽ���G$Q
m��1���w{�SN��G�z��|G/lX����E�ۡ`Ջ���
��9˧>��4j�J�'RnR|7UK��B)Tb�Eu׬�9��Ѯ̻��6g3q6��0����n0�S��AX!S��#�{�C4d�45����(&ʫ�A�L u�A�7Z�%_�E��a	$<@4EyN���tP�m��M�`ӈ�oUisX"=X�$�����j�6Ol� �%X�� ���r�d?��o��VP�LO�[�y?��
5�����T'���Wec�tt�9��g#=ӹ�JI��p�3|=G�}+��l�W]|����XlxVHYEB    95d3    18d0w��$�D�VzGd�?�a�dCڕs�{� ����9�Ț�~@%��V�y��� ���(��[aB��qq5��6��^ݜ�rp��T�W`�>������\!b�w�6:�����dC���QH�Zޞ>Ȩ7ѫ�Y���#}��ǈ��(h%����O5� 0�/����T�G��oK,�U���GB��5NẒ=���96�����3��Z���t[s�
����������ޔ 滪���z�Q!XII��L�����b�i��v��)��;'��{ɸ��X-G\�Y[�����.EdX�!�P�Eu<6�d�"�X��ǲ='�����){���:�	�]
�O4�i�y�e�Dg0*������-�����Zw7�;V����I&�}�K ��k�ô�]��,�}����Ү$G�u�	���E��qeظL�B/٥����d-;�n��'LU$�z<��ҷ0�b�Q��O�����42I�E�0~�>jE���pT6�E���}��|Uxu��2*�q�x��> �\G��\R~�+������+�%�/�$��늢W�p��(��	�EѰ{��\c�P����=X7X�n\���[ ����t����_0��@�u$H�]%Ԝ������UQF��.{/�4��n�_f��lW��f���%�!i�G1?����^�CYM	�r�*�}�ܻ>�n@����=���v'!�h �fz^,��E;?����Xt��?=?-F׆I�qY����������67����9)�>5�
{ᦑ� ��!cxN�b/�L��&%���x�:@�������1*�����s0z� :�y#uj]^;�h*A�KM^g����E
$
���#Yp�U��v#&��4�F���!��zb�j"����kX
�H���/0R�)��ݬ�z��x�S��̛�0��)�� ���x���k1OL�9�4�����ͦ��`���������0F���&6Pg1Bt;�x�~{��!�\�O4�+����#��ҵT�T?�\5(a��������.�b:�#;����[p*l��L��S?>�%�'�iP�E��^,�%�-�A�B�LY̿R�!c��P����0�C� 'z���H[1Qd����kí�Tpdt�D¢&�^�S���_i:�E��&1�ҋu����2�e��`1����J�z�1��Kjݨ�W���`�X�l<���y̯n
.�a68��r��6�}�U� �cAV �ȷ�g�y�u|�7p��O0�k��?Z��b��֞+ws�V�=Q�, ���򤤒5������Z���G��@�A_.�-n���=��)����e8�a1�*HŚ��+������N:�`���T�ϖ5�a�&$��#�ڸ��!�Jr�_�`�)�W��O P�E��H���	��-v��u	�c�5�4�g_Wrn߃��Φ�z�	1]�Q
��"���aYk�J�Ag���L�*mu�~���E�R�}H�%�e�;�`�D0�ߍ�xnb���8yn��i�C�dhx�{xB�,�m��f>�^E��ܫ9�E��%��wVY����_�"���D��Os�������I�Uo��vS1�"�-3�O����/pXΚ���Z-e_Wa�E�OLV����Y�b\+�jcC����Y�H� 	�
�H�Q$g'���j8�jRc�%�z!�TV}��#�S���?������6�@�D��Jn*��O�f�U��)c:*�7o�o��؛�,���:`�dn֒���;F����W^.V�D�HM��V�O���r��؋�F�9w@H�0@��㾗h���,�2E��9/_oQ��E�(D���Kh��2����SQ��i4�M�.�L���{�K~yP(�E(^ͳw�'.^p"��K<���
���޸t�]���N2��i��uK���{sҬ޽da�[5r
�1��M��h=�N�]�$���32��'��r��$;�/�|72d��z)����RM0s���E���1���������6���k��P���y�$��3q:e{��d��}���@��j�0YD��WV�V$ՠ��0�GNw�Pp�4���٧ȋ�A�|�㷚R�T�fĢ�_ D'�^�f��S��2d��AV�>����b�;Z��'�S󑯄�b�#I�	��]��OPA���$�\N�&r�g�iV�A$d��Y�����#m�T�4��&�|�3eX���z���$���J6w�%<cs��|�]q�3�y����\��/Gю�� �q�7��Ҙ�N�u1>��f�_n
җ\e]�u�Ҋ�o�W�t�Sxm���&�6���o�C�j�{�,���(�(x���Bl)�D���o`�P�«��E�ٹ���i���ں<�d��	���j1���;�T]rP�[��e�%^�(s�im�E�)2e�N�1�b�_M&!��Z�JK(2W���Wt���A�G�t�c"�~��?f�ٚ�h6����5y6���=�_���,/�c��M�و���0�	��FT�?����龷����&2%��n['P���_��	�B8�Q}ɀN�>@��8H��x�&?[�p�����|[~�m�\)#�����S��0@�d�# ��C��\�����[�>���=�-Xɭϯ�2E�h;1?�q���_��lbک�=Sy4S>P��y�(�14�z�9CU����m�!����%��C�s	��Q�,׼����·&�Zנ5����L*bN�����)������~��$��{~5v��\��
���*��Jfb��s�,5�??7��Хk?S��ޕ��8�S�?�em���ԇaj�?����BY]���Y�E�(F|��>���4#�o���锢�����)�x:@�ڛP���ɄR��dQӲF�,�̻e��%�ҿ�l���AI��s=���~u�����q��m�����XP���H܄O_�z��? 2�k�{JU�a����JI�_���)WW5�¨p{!Hj�Z��]�!4RR 2�����"p",wK"q��(I�5s��g�F�h�iu����Ysb��rgj8�X�:�9{�ZW��L�vF9'�I$�!z�H���3Ʋ���E�u�O�ׅ��=O��=8��M,@h��!����})����EM���m�93N+@�<zӞ!�I�ө�R,��|��ߠ�ke��(�0N�l�3���* �_�Pr Tz���������i���E�_�x�W���Φ�����ck��@�O��,k��AF��@皞{�`-ɑ�u��x�<n��T�*�~�X� `6m��0ua*@�1��[�U�H��0^�
�[�2N�G�,��vb�v���diP=��iHB�q!�;mQ%�����u? ���1x!R�_DG��kg(����0UU��P�3�ȉI���,��Jh]lB���x�K]DBx�H0��xM�Q��eޔ&zD��/��8�uJ'уnFu�$���~��茋~��@-��8P;2A�%�d&��p�t)�&^k1|���B��/� �U¼�� �e,�M��	T}�%��Ĵ���Λ���ڶ6�����Id�6T8�d* Քn4�┳��Rő���ͭ�6m�L[�9� ,#��hX��p?`;k�$<j�^�6I4���ަy��l�P�\h�#>�D�iPy�>�K$K�.-��`�$����ӳN��pp�zU���	�>p���w�mx$���,���鄅��ٟ�*?	^%�J����=��q�X�ȓ&I���ѧM�İ�7�h>�Ҵ�lg�_je�޶^�2�H׵���ZrW����BYrI���������V�x 6��(�|T�O�B�h�G�XTh�t�6��:9o�UE��`�_�"�+��e��~oח�V��S�2&V��U-�!
3O����G���/�0����i�(�?���_e	њrH���x���n�Q/��\ɚ�;�U��ߋj��&�rP��^#Jb��WL��@�7ĘZ�T�1}�4F5���� cd�:g'||R*կ.Z����R���o\9��	�)���(�m��T0��G�J�Ulk�D��t��J�r04z�(�Mx:��#���.?�W�}�$�}*N1��������T�@E������nn��}ח:�{%#H�1N��xx���DfB�2����F����>�����L��n���9�|��~8�ܓ}���A�!(J_;�M�J��,Wb�_�T���%���k�D�I�{L��W�����^!�߀o��!�P��_�υ:�צ�V۶0���9�\����'���+�O���m�ZP����i���_�Of��^�N��w�?���\6d9��ƌ��V��׾��q��󺈑"�3��ǥ`H�$�1�rr���qƿ�y��&�)y��p>J������h�Ũ��-�����x_�����G�U}j�����1�����_Q��"+<"/i�m�����7��֨趱k��V�N�]1��q0�㋉��d%$|�t��n&������KH%{�Ag5��8J�f���Xo[�l�W����be�h�۞k�j��%� ��<3���57mU;�v�����v�']�d�[�P�J+�v�Os�jt?�'�hv.���z]c��Il���G�9�6�O�u@ZU0Wz��$�����hg�9�W��\f���3�'�(a���$�PŉY�K
y�����yX�����Ou����E��9[&�P��}T�)�o����S�`� 􌇮d���I��q7-���Tq�|��;lh�
�\� ^L��U�7�>�K�Pా
��I�-�`ґ�'�h7�W?#MD5��ڙ���p/ב��wUΣ�V�/��7�L^]���*Z���Ʊ�(��)X�<�~I��:Q�,tu�Y���_��8Y3"�-&���X��
��0g3�˳M�Z���LM�Hƀ��5�$�i�i��g���'���k��E*i}Uq���XuQ��G����Pm�N�����`����=�Xbw����#tֹ��y��2��G�6#UF���v���p��nır��7;��t���q.���c3`�@q�3
wL��D��f�9a)��G[��X
?B�>�X�e��aC�n�d����p��]۟�F�����ܰ`�ez�P�F�����M\�x��O��0f�~´{%�151�$�I�<اw��<>ω&��+E&t���ݛ�E磊���A|
�l�{�dx�9��XȚT�����k�i@��]a���`Y�4�?(�W�m��﷍����3G�5�~N��qu�Ųƹ�^�r�_���h'r�����mA{0_��".'��ޏ��փ�pg.7�%�B��5��݃��2&���o��;lbBI@^�0@	}2��1[����D����P]8��ia��Б��{X١���2�v� �datc����C��f�1��fG�w�%��Ks2�FJ�U<���,�)˳J�����'v�Mg��1�<787�3�oy�=5
(�(Ų��kv�����ru:o���7~��9f�R�������A��߹�c�M�>����	���ǺF����j~�ͣN��̪���*g~Q�Ii�?�V�T~��H�Fd�/L���4��*4&3���L_b)D���-s8N鹕 �|6+���w^��R5n�/����'aM(��!Ʀ�I"�x��*F��q��ݖװ��Xv�e�nA�m��<��╗���V��v�I,v�w�#@ �Z/���sb�  �f^v@C_���-�|���;L�����AA�ế��hZ��a��=S	�}dwl"��.���ywY7Kz_��̼���
?SK ��ts�"s�\�Zꀵe$@1��m��bDv���5��޲>3�pԤ
�&b�;�8�qb�Y�2r7�ǑX>mt�\p�.�O���i7�����Y�F �-������L�~���n�&],��I_O�\&$ѥ�{��q�T�乱����rd��}�[���Hs]4f�y(�h3���
���[&H�^�ư��ξc�xn��5?���=0^�(��TXG��7� ��(I&�rS���"c=\�#W�.�P����#u�H�p@��ϠE�S�"��[�2�ݗ4-��t?+K�J� j�I�~]!5�eǙ�6]R�4��b6W��X�>�>*B�\}�(��޻E@�y��p�'�#Y0�D�����P}7×D���P�H�_O�%�J��