XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����u�ipt�,�0��g'��ʖ�,~�#���!��>%��`Vz���ɤD��Hϒk8�]����rsd����x��Ϫ9tM�\�f���<F-5�@ّ����mc����]h��Iea��\,���k����2�v�.uA�'z�.��o�y�.lM��du�o�t͕��`�½��W?[֕rfG�Zez1��aZ�r[X`��:Q�I۾o��?6*{*ߛj�9
�xU���Ű�����r{s�
��uT���zBe��>�5Ɂ�����D}E�[F��Wn����J�x� R[ňL*�:gI$���T踐n����#�[�����氇R�M�4��5ށ�{M��-	�����D�}Ɗ�k	���O�W!ui�X��؀�)���$<A�P��ĿF�g��o��-���� aa'20*q[x�����cY!��4j��8�g�kT�8X��	�!��;�����>�an�}���U 98Dl�ŀ�2Q�]^�v*G�D*�z6���SI���+OY����5w7U����� ���O{�_w��cx��~Heb=9�S=�^$#����Bx��U@��g	�:�u��Z�:�Ӕ�V���~e�Y�hE�!Wj!8�s����~3]ς~�	�Ƙ�ET�#��"�ue
��U�ğ��䋆���,�a;�]%<���u\�&eP[0F��'�E'y?�t�C��ܼ�bڑ�X��1�/dg�x���Hۧ�)�%�ü� �D?��p��:��@Ʉ�[�XlxVHYEB    3e93    10b0�0q��!d�҇�j-N�w��'��j�����5Y��:�1���Ds���r�LC�Vp�P��Xˋ+����f=A�W�d��gq��_g���3�lV2�Q��/����^C�b�;�W���n�$$��;�'�Q~�jW��E�d�!+U_H�J"J� =�r�간��̇���!���/d����^�������aF��G��i�5�6KZ�f��q��߷���ce�3Ãp��ͻ���V����x�D��9�Z������[�fdo�u k�v��b5�VT��^� ��G�>]u:�d��e��ώ�����V ��(�O<*}��t��&W���sr�U���j&-����;7�?�s��e�47�%�:�5�
�������M�|�hV�8����b,g{.f#Ysȍخ�,�Y������)�m�ڠ�k�/��j#td��t�9��(�)�t��}p���I�1K�{�I\���װ��Ï˞��
�{YO-�_�
��N���I��ǸKZ!<�X_n��� ���JH�!FO��R߭�}59�	+�Ã'���Y�&A�#B"�l����cM~`��u7�h@�LJ�ۃ
�����q�Vi��i+I�Gy�!ae`�D�0�sc��d�w�K,�������/�>��"6��0�T�/������.���n%�>�ޔ`��*���[����[�
�uW��z��ُB2}��w���7fsB�͆��~�(�6��Pp�D	2jY8l��7��
�%K��x3
^��;~=�2F��]Je1i�UM�f��Yn�W��<rQi���I�D_�@�������ږܮ赔?�W���Tf+�=;��Zg���#�qIWyyW��Wt@s��j;�s�W1Q��0�
��#CF�1ѐ�eel��I����BO��t�,ӟ��p� *7BE��	,�^
�S�Ӷ0�tR��
Gas��0,�t$j��g0>�L�PT�n������v��4Hyl�B�c� �|�g�"f�A�;�]-g᜜�S�ߣ��B���;����ϥ��g��D�Q���4�`yK�,>��v3��Z�m�uC�9_���v��?$�f��y���i�ɬ�c��!;SU<otF�ḽV����b�3|M��1���wMMr�O�Bw����L�Vd����c�=[!u�(g�>�	B����(�^��!�� �U*�`���BW�:GDcmi��/��p|u��F:�㾔Mj����"�fm�?^�Lg;sŃ�k�Ru�9��� ��5T�X�	�#_���m�Խ=�[��B�������)�Z�gi���@3ͦ����|^0q*�&�͆�1��������lH~2v/�T8�o���V�y���Ԟ�ā�s}]ˤ�A�60�D0o`P�T��M���ag��ge�o�W�d��!�Z~�}Y_(W�e�
�#r43�Ó�<Y�[�srڙz�α�F.�z�w.*[#��X"� �r��X�Dd7���k3�(��D��ʄ����nS�y�`917��P��HYO���aJM�B�E�G- a,���p�.����4�dB�/�A�ڨ���ʮ�9����p,_��<m"_�����o\���BE]��]�h̚�74�80^T�G��_��!���ak�A���.��	đ�����t�*�����mdv�.��c�;E٩J�}�ؑj��,`%N�՟�}{J]��7W�I賠*ˁ�0H�TCm��ݚ��_�}���i/�Vo;�:�.��\j�|�)5x�r��9�[� 7/1���U��K�߭���a�EX�t�wR�o����Nn���=�2h&|0)��D����#���?,��Q@��S��rYr�������F
@�s[�K�^�"|�G�l[����v�4�J.�M���3:q�L
V��p{F��8Y��(�,k�6��%e��l��z�cе�����<a�@<���Ʒ��:�w�%DSkS��� ��gθ��R�/òr�Yz��5z���+���ٷK
9���/I��e��c92��`:����ĝ�[	����z�2���O��آa�p!��^�W�ӱ��kI��^���W�w�3*R���sµ�?�~^f����ץ��U�$��g̡���D�z����	0������'.d�r{P9!V�]k�����%����v��/nb�ͦ |�Z7ߥ�5���yF<_�/y֊�˷F_�?���V����Ⱥ&!bb�r�F=׼������1�����ȹ�g�6�0Ǖ�p%� ��;W��(�����Cҡ�&1��jgP��H�m��������������/��i��M��j�!�\�Հ��,;Hٵ`�������-�VpE�*�����&O~vDOkv^�u��ML�֤��)q�E��
���,�ő�"�0dbHZ#�0��=�V,A/�P�O�� 1�'n�KE��z)Y�H��#���t�5����@�L���IP�~�g}f��
0Y	��h��H�|g�Q��*=�R��K?��?ƍ�v��u~Ì3]9H��O��ϝc&1`HmL��i��3�>u�W7l6�E��I�c�D��Hs.k�Ɖ�e�L\��z
K�r`��Hy�L|b�ڎ����.�L;�ceS9���8�����6�p�F�894�@�4+�ۓ����ĵ����s������lK��!��D	7^��蚙S���괽�A�	���ČLD�u��a?i�:�<����c.��Iv�����P̥�L*_���>�z���/�WA�LqM�d���|���1�!#������
b&r�W}�bH�%���Ԑ	�qu���Ƞ�������%�
 ZLO�^�N���y�,W���̪�y>v�c]��qBZ���j�#bCx�	_x:�ӹ��bC_N�����	.�*�L1GX�:�0D���oU��v��[Țy����Wq�^{��m�D�B����1�^<�">d�FM�l����\/���ݯ��x/e�f����j5���y���y�7��WQ�Yh��?L�Q�	l+�b�f���2��ׇ��o�X=RX������Тd��ȽB�U�W�~�Y��uM05�T�`p�=L��8�WRW[u�<�+�[�Rm2�0Z��er�}�*o��R�as���R@��.��<3W�V�S�6q����]p�`�rW ɇ>Ή�&Y�|木¦oN
h�C�߃��hcHT�쒐��ˣ�@���~$\K��FwP���Q:��QЙ�ž���BoU{�"l��K^�Kc��אA1pmr|/=��A=����H�Z���ۏ[�C��-Ћ�X�h�
,�2����jX�<q>���qj�Z�B��f���e�A���
��S/r��"�,�"�%2�=�	�>%cj	�v�9ٟ!G���+B�|Ů"v�b/XȪq}Z+D��ۚ<9�Л��҆�ʇ]���҈8kb1�_
d
�������_��J�{4���0o}k�мA���t�	��0�����%h+�[��A���f���r�o��B����Ko� ��M���ތ@�3Z����m�W��ebg0���W�0�O\��,-�g��T�lnlع~���!Q;�w{��E`]k#~#�"�|65l�wjC@pQ雩�^�Q�L�~Ӱ"����i_�*"��ݏHQ1�hd��>f�9	\è�E<KN��>��߀�o���a����}�Ď�-y���Y��6 XD��=Tg��`����F�x��ǣb�7�ڠ��w5®��h�U�#=�����`�)�I��UY_�A2�7b�6�ғ�O\����ϱ�J���z�U���W��Ҿ�[O� �A��:^&WA�@�����fI���i@
��!،+�����[x�u5(>���U�Қޙ�_�$/�O�ɫ7��ݔ�
����ګ�`Mm�Zhz++�wQ���M>����\�����ï
`r�.:�%�4�u��?�զ�\��qb�AF���Yu�t\K�����%����7�yR��7#��l^N���L��~=���P�/���+���>���ϡC2�7�v��lĔ|A=;M��ޤw���Is0��0�PF1�	�/��);�I�XC�Yy����I����<�1M�}�I6L��B��<W�$Ej�.Y�;]�RvG�0���,	��k�#g/AW�����ֽc�)~�I(*+��'��B("���s	��Cb��)kʍ�\`�2{T01�