XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���[�fp)����0+4�ݕ����_�q���P�s~j�_z��62^E���N=�K��+��X�]�y�q�1����ь��*m�	�#*i\�B� S�i��pkm덢�l̵���K��W Ore�E2_ؾ>)O��2(�/��cuo����e��ЎD}�B�����W"��i:E�K?0���E�E�0H���2�h�|��ȓ1���D�����]Z���=�	^� ��P�.��-������÷T��a���n-�b�Uՙ��[�)g �gr����q��A����d �qE{�ӈ�+���l�W�5��
W���o[y�e��<�$3yͥ_3��}�>[\m���
U�L��%z�z���P�3�yrԳ�\��vn'X������3}F��R�����,��{4p���]�J�jĆ�$���:.���*��*r ��P$�'�x\�D!,x��se��R�-��6������}�L�i���5��U��a��r�aG�"A�,٩�6/�I�0(�S�+Q�� ;eG��`��1��Cl� �ŬH�2=�t�LC%�X������A���ԐJ��8��.�4]�����τ���h�{��r�rv������de�	Ie��<z;�4b��D��VOv�;7���e��IƘ�Ki�����ne�"SD#L��1�c�L�5����%��%� �g�a���T����ޯ]�)��8[�S�wad�3�>P��1�sZ��F�Ź����%;XlxVHYEB    1448     800�QMXT�2��H�>m�&FE�w��ıvZ� �G��ߘ��5 �f��Yw�޶���4��;<�&���j�+�T4��҄ź�@-��zi��ݕ3Lw�#E�<��} uM'o�SJ�Cɋ��yv�E������b���z��3xeQ�:�f�r�#�]^g0/��k�u�P��Kt�U��䶑t�q\��������\�1E�	�d����䰆��6	c��f�fS79���~Ƈ�0#����R0?�����pX�����:������K������Tk,F�G`�U���D�k��}�ԃW�`DL�<.��/G���u���Gf0�~�2UA1L�C��@���,�=�%V����?/�{��kr(k�^�`��x8$��L����T�玷�yʑP���@�~���Et�D��N;�J �-����b&w5E0{�n��B��+�}�^���j�yO�<��`D�.��6
�>��O����~<X�X�P=�T�l�Fz�)}t�\#�_4$����o!�b1l���(�����`Nn�ͳ���ǐrhwt���I�=���Y�m��HہZ�@�ut�dk�1�"DY�l'E�Q��^'�i@x�,�b�!�רχ�))�����q!bj�#�N YN�p��_ت�s�m|0��[�w��O��Z�hTy!��=�Gㅙz`��	ټ�(]a�|X�=��m�
{b�@Q��م�!L���� [V*>��l��%h�?�{u�������Q�X`5w"ׯ�h���?�_I gj�~P�n�r6�Z�\����g�3�zΓU(���Į���>���MU�C��.�be�����@�g��l���')�;�?;(`���#��U_�Z�u���̄P�����1{�)��㘜���z�l����7�OY�0peK�I�k��9	@��(����@,�W沝���dVL-#�E��Uuw��B[>�ϒ=�I�o��	��o�'t��u��3Ꮖ���m(��������z����?p�-������A��5>�4���L�7�@�����F�#47��y����U�n��`FkQ0<�OK��͆�ը�A�Hš��7��j�ღM)�WLAXg Ү_]��-��Ȗ�����ͦ4��1��"�4���.%a��1���xZ��4��T,�:��#ǽ�Ǭ]-"#���:�B��ҫ
���=���!9��j�\G�8�Bp�>L� ��X��ae�-�e:�?"�dF��2�c���ѫ��	ji�=� 1�xid	�*Dڱ�_R���;ؠ�����Į�s��q��h8�fѤ˝�Q��K\��h1�h��V�}�4���槏h�/���Ë�-'���n2Y�bb:��eN��3��+��D�aU�ƀ����B�q��=�H��¢�a���L_gC��_9�X�7��12���@���/�0[�*�l3g���+�<�9����d�O�d�y��D'��cT.���WD� �R��g4 .�B]=��d��l������ �:��1]�=��ˢv^�hv{7��gad�E���S���Ա�p�Bf1��p9?!�!�W�O��\��tOQv��bP��%��{��.��x�^=ק���3I�bX��:�A��nG4b/��P0AOh�񕥌���6�7�`�'�����n�%]N�&�n��*�Cǆm���7tDbx�� ��X�.��!<�gKل�$! �~%*
�Ż!���Hq&� <6"ꥡ28j����lP�ʐ��N�!�+�ՋE�	� ��?HX��]�,��<F �H^h�z`��c�d��4��h�'v�pLS��BG%ͨ`b '��ui_��, (d�SG)v�gBQ��"��Ok[JǪ���W�W��k�n�{[��D݃7�8��^E=�w�s�A�w�~��7��tG3�tc���]��v��@���]���޿g������#�A<׈�±�����nV3�2O�Ċb�}���e����!�Y?}[�Z. 3���P�x�I��#}��
��S