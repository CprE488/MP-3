XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���?��:C�VjJ�ف��e��A#v���.��i�E�M+�|W�z\���}��z�G�����]B;�l<n���ĩ�׿�V+�N����^.�>�J�l��|S{��ӻ�
����K�FL_u]�n�V·����J0:?z�f0�3�m���S���|Nl�&+6-���!�_�pܥ]��b�:���"C��KE'�2�Y�}�E�%7:kv��+	�����3�>(mF�����.���DR�%�Q}[?j!�z[J*]�m��ҭ~$�''\�b�=�Ѻ�N����F)��Y*0NM�7�T	���&��wŒm�Se<�����ƌ�';b&{͛�q�l�?#���T���k��RM���9땒��Q�?fx�Gt�����zE�@��&x��}ę���g����8�y�k�9�{���y6B���io]���ޕ�UQ�.��+��x�-���R3/$�C��:ʒ0'/=zQbhQ
�k�®3>��6]����3slv���U���6B��i������u}ٵx4|󩺏����2;pT�,z��F(�Ԯ��f�{j���
^'�6@�F}<�v=��TCLk�^�>.��No%s4w�cM}h9o�t�y"5�=;�3L� /��>����y�f���^�S��NU���a~��i�� Cy���LO�"~���:�o�/h�\��������t�w�����^��\c�h��0�ll
"�N
�C��Pv���G��T�Y�����+5z��<x���6��bXlxVHYEB    15b2     890C�*��_�>\&���Z"P��	7+��^.���	6�m߄@N�)�ݿ�9p�W� �&�s<y1�������%b˯ �����Q���|5C��oXߞϬ:�v��Y�Fi���u����x��ѱ�N-�5KR�BA&F[ɏ���(o�h�̤Q���o�K��N�ãP)5L�eo��,�-U��O�y\ٚ�$��aT����+rvl�~<U��T�k�ҋ��}k�`5R#�U䄹$"�_t�Is�?�*,q��6�q���[�bDw�Z������K�t]�'B6��\�N�>��nְ:�{��T�-.O���i�R�7���p���Y.��-���]��?��e)ؼ�������3nƏb��Gv�j��y��/�hiX��5Y��I��D0�m�Jz ���R;����z]��Sv6�F��8$J����*�����\_�#��%��
�ʳ�D?��7�J�I
� ѼH�%�YD1��b��*Fc��eF.�
A 5N��9���A��927�)e�ڦ�S$V\��������Ѫ}U��/͖V��Ȥn�eQ���\��}?��=��M6�e?7]ԴR�=:�w����F6�8AX���g���z
�B�����?3<�}�s�"ň���/�/�Ew��Ǐ+�F?
��C��\��&E�k<�%�{��~���m��9e�]�I~B���*�q9�Zm���� ���g�eT�3.ʝ�]���ŭ�Lb�ś�*�h��z�����%i�A95)�s0�G ���z�m�
H�ۡ�Ͻ��"!<�sCK7�zχ_6�~�O��q�����ל�1�?� ��u+�!��so]�`1v�:���5;�;��֣H���o��5֧}�i}�#��
L��ok�PVv�LcS�daC����!K��G����ݿԘ
��=I_x�F�@�,�CP"�C�03���YMl�u��@!gH�fJ��J���q�.$;��Nܨ��ޜ��L���}��8���$�����a�*^�q��M"���}:�]N��0�>4��O��~�,�����H�2�gK#/�Յ}#��2Gp$˙}e=�MK_g�����Y������c�B��ޭ2����mFc��w��X0�������5�T��o��As*��)$H��zKk�ר_�{
�|�a*�v
��(ͽ�KWf<l�Ǧ&�A�P^��$Lێ�~�<�H�R�3M�݈u�a:���W�v
��?�a��[��D�F;�$ˉ<)Vr�E:.�Xs�v�.߮�N���J+Ǳ
��ܞ��|}d�t^VZh�kN8����3�8���F<3r�~�W�c%d�)Ag^|�;A��C�?��|���1U1�6�(�h7��
+VjI�K�_�+ϏZd�uT���E�jT+�����Hjsy��p�9-n�U��}�{&����0`���ӂ�Ɛ5s ����f�~�і�_z@��[G9l����~;#4iGNqL-�a�G��cy���w\��G�>σFE�A��)v
,��	������3���Q�D�UE�x�noh{��0{����C,țM��B�-p���]�[P����Ԅ�@
ˮ�,_*�*oϛ��u_���0�	b�y��F���Bn��qO�w���>X��_��R��ϭ��gq�a�v}�#H��SN@El�g��+�o^�6<��k���A�Kz`�`^^E�����A��s�Jp�5�Ҵpy{+�A��*;悘2�wO�c;�mґ���h5+�ӣ�[΋C��^��e�3ƋJAx�Y�� �s�:g�\r�o�C��e7���:V�F��겂-��é{�ª
����a��#~�˹��F�tAu��Oޚ��,Vqe�C2W��7f������g�*J�&�6��&� /�3���8�Ms�,���ܫM�ǖ���mٳ��=b�Oס ._�s���Cu,�Vh����x<}t�JC^Q1-D��ώ�MQ�A��Ģ�(Ś��A��
R8��,���M��Fb�x7#�!��uK�ka&nd�?�Ah�7��4Ȍ�{X���Gu�߯�&�zr8 Y�q}�c�sO�=0�Q&��}9�(G��aY83�J��"9�+Q�Q~y\G)��~�����<P~a�7��� /mrɚľ5%��$u,��´!vCX�_�3�-�%�j�N��дĚY�\�