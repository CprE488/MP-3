XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���%y�#R�k��YoX�m��кͅ��Dj{�����B:h�х��l��P����T�׊>�X�w��5���^���k���W$?>ߟ��akg[�4_�r��D[ީs�p�j���wo�����ϘX�����Au-��`�7=+��b����>�T��`l�7=�܆�I<������d����\j7BD��.Z�e�b�L7�&>L3y�Hf��h�-1�3�<�m���6Y�!L�ЙO
�������%# ��p�^ n��h��]_}��}�[���E-C������q�<��75EF�>��؍��6����֙6�bX�=O��/೥S�=��(0�S=<N��?�<�l?( �nS��<��m��.�A}#u̐�Fl@���S<��	ݿ�^��\�8D�-U ePon�Į��Y�����tI���c�X- Rh)�u�R�D��ȕ�e~v���U�<�.���[���
*WO�ߟ$˺�P8g�䣕e]��"�b:+9�x��\��7�v�ÉN��:�L������a�Pv1�x��#�`��d;8p^5�J��k��.��v��:�E�����5%3%���	5�����/o˒���4�(�1N��%}q����I�3����D5Y҂��0��d�A��M3wB\�џ��Q��2hϮ��]g�R��f\~��R�gY�*B��3R��>¿D�j��|�'�R�a�gG���|x�Gڬ���G}!���r��OX���ø�g��R�I�~pm#�XlxVHYEB    82c3    1970C%2�DΏ,��;i�qU��|����H�R�Z<`�I:��M�R�!�E��aTc,�8A��w7��Y52�Q�}x�[(��[ܲ�*m�S�o�))B=�*!�cY���SZ�$o^�@�@`w+7��"��5�����W�yv��������DE)����z�_�x+�p'� �����
�JI~H ��
�Z���e~���xx�Lm�P�']6�����M��>��%���l�c£�"~�;;$�;����M4"½�ro|$<��I] ���^��x��jF�,��zH�!��Y<�ط�kM�B�7� �y�h�z �"I!n"��T��e�<"�I<�>�d_�I��cĽ���ƍ+q_��.$.ׯ��9Ļ���I�@���O���SYٸ	��o��r�n`��p���N
�����upݕ.���EˣRP��4�2nJ���&�3%t��{�ZN���E��8��YN�e��D�x��7F��(�k
o�4�;?��fU�V_~�Do�(�%���R�Jћ��f��^�6�K�D{���"g�^��*O
�׵�I�ƢXoZ;-�����ǭE��WY!�H8����2?D"����:][�w:>�_h�z��Dc�yx�ځVj'�{��m� �^7�*�6��دt��Ɠ/�Oj����S!o�+���
�Q����1�����2��%�D]�S�-�Q$��_/��K��f��9,<c�S��#I(�~����*���;������'-.T�9���"(P��Ճ�8S >qX��ے��|��<�\l�xy����)w�LW%�?������D{zD�eV�ݛ%����sMT : �a۫�e�|6j���c4���;�����;_�o�J�����7�� p��rN��v<={������a/W���@{�8�ǐ�n�Ic%�/���A_�^��=u���}f-#1Ӵ��m}�4O�0��0@�n��e��"��?Р�����IM�wԞ�sz�X������þ&F}	�Li�dn��l��r?�S��i�1YE-Y�Ҽ�Zn- 4�x\�ak#�?JI@���^��|\�J�#i��&x�ޑ
��1��U�aU(�ĭ��nm|�/sݼ%[�*�������-O������m�k3���K>f[��TE�%��/݌/Q���v�)c�g���7�䝍SwQS�1tK�yIfP ��X�+g���5�xbX���5�C����WG��YMr1*_���zB�v���C\
d��u�<��b���"|ۄl�u�t��q_�N�a�>�΋,[w^�Q��s`/!k>�j��Y�룊L<Ċ�/1M��pn�icK��M}`��@�2��Rq��rṟFn���toa�o���:��>V�fob�X{���۸�N��M���>T~��l�o�D�lM�B)�Q�����<�)]}zUF���p�6IA��>&���Ǆ�KO��$Y��l�
%��[��΁�����c7��1���PЩ��	�j�����?�Rן�=��罴GU��8�'��ޖ��R-婊��4�B�u֔�~�H����L������O��1`(�:�EN���d�����o�ҕ��E[U��w�#�1���9\�&A��^�������Q)���M�]|�/�ۦ�	{]k���~�� 9�o��%�ה��$	��yj�W����r�I|w���G�zS{���ש�����t���V�'�č$IC�%O��P�ȴ^�"�� Tn�[�
͒a��t�a�b�IA�U��j�.k�+,�d�d�@k�7�k�L5Nz^� f	����Y�=�<Vtq7d=Ϭ?,���@C���dʷ̶�WWݵ�uU��U{�9M���d`��n�ˈ�����2"�~� U�H�Q3��W�dTPmZ��*��������%V�%��'9�%ߒ��vs΀��9�/�B�/�-%v�\j�ISԽ�;��%E	LЊmO�o�4�y٧7q\�(��B��c74+�X�9�������!�B�Ë����@����جòr�^
Օ� �Vv�ım���R��^8�Ŵ5ޕ�(q6�$n�1+w�7�P�~&*���r}J��6�~��ؤ�w�@�ߞ��QM[s}	a�_��\w\	$��q��}7������Tq��Y@��y��f�oZ�֗?`A���+��� $�����le�S���
-��a�k�P����r�q냨��Q&�砋+�h� ﲨ��	##�Ol��g��~vS�gJ�Z?!B���������6���G�NpE��г��x�J%�/�����u�CpN�z��8_0�xT�Z{dy�.�d8-�E�> �p������g~i�$]{��F���V:j�Z|�	��#W����-�b��l����T3��tS�	���67eP�G�d�%9���
�/M4�"�3)��G�N5��Ч��\{�B?18"��i��4/�2	p��ے�M`��i�sd7�6��][�we �8�;)O9 I��J�&,�Y;���]P�z1�߲�:#.|����%���g�����>�N��#L�I�c{��+�� ,�A��ȮWj��L'e������h)�|Y:��˺�=2��걇�8�������F	��6�9��uLXP��N�'cI|�/)�#�y�M�=��ɑ�X{��s�9��g4յ��#7/F��)��_X�z<E�
=���K@�]L��]JA�}z"gKO;����?�/���&Ͽ�kH���-�b|n�TP�^\س�}��8�`uA�3�mu�:�W�k)V�-�&7�����0ǳk�L�98���U0�wW����3;N���7�ftV�\��1�E�
"��@L��u@Wt��&>w�%����k�KWR,���p��^��<E��G������[ :�:���壳�����q����8��a�w��xF����.�y�M����߼�Q���5�� ���at�~�`�hl��4;�PYдA7ݺ�"B���
�Z��d�u��B�Ё��MzIn���b��M�Y ��7޽�t�
"~�	��<�n��I�yAųgw�A�/w���˶���tl�>`�����1���C�"/h{�T��7!J�[�M];��|��ge���K��\nJgݢ�jv�+��A��f���*���6KD�~B���YhݘK�.G�e��yqI��Q}x*�i���:��Vn}[�|[��J ő��,�U)��Ҋ�=&� y�h_�Wf�N��S������Ǔ#G����b#% 9�A�&T�����4FB�J6�}x%Oζ��X�g��\�$�9�S��v��������Yp� �Y��뽯Ry�4F{�x\�� I�īRqrvPlC���J'�?ٝ ����%�)Dqҭ#v���㳃w�e���E�a��f�<w^������ߎ��7?��4���As� !�)ͥ�a��E,�|��k^1܋jT<�`%��Pn��A�r_�����Q^�+�zj�|�m܆9q_�����=����&V��V�����¡%��C3(~����7�X�9�De��'Qg��p,�b��306Lln��M[}�}�����6�z<���&��)8م>�5`>f<��L����{+Fw��~&�P��V쐶�[�r'͝��M���U�l�
Y������b\jpl���j�iR4Ԑa��Sۃ��>h�.� ���ř�ŝ�[	�B��ӹ�KM�ܥ�F��pV,{�;-��\N`�n�[.����1�*n�0�^K.-y-�ze	rڭ��e��q1%+OfkE\gLA�0�fX�����?e�&{�A�����k�]'��d3dӓ]0z����2���I|gk$��M��s
�����tDŻL���-��rS0ln B5�ɞ"�)�a��j-e�oz�����lc
���V>����V���)g�;�|�/7�4�A�\���@��X8��l2˄��8�J�s����Bb�HΖ��=�bK��m,e�ms����K�*j���8�u�}�j� Î�T�PX��������� ��X�r�`e������=I_�r7.'�6*��D5�Y}�YY�w�.w�ZZK�PkJ: L��Bܿ/Դ蜊��6��n���+1�Rk�N-�m��)�b90p�Ķ�\'��?S���S/�#c��$)��b��j�vy�-o�7�w��u ��Ols���nszg��k�e�a�9C��WU�H���R]����["���9�t�@\��D���40�",vYj�x��>�"i�JY�g���`14�2�r�(�:q>�7�7;�.���#'{	u���i=o�d˴�~�M RQÔ�u����x�N�C��hOEY�ـ�l�<B�>���9�S/��uu&5��r�����H,8�.���H�|�xR�ґ�nT���>�1WW4Z�zޚ�_��4x�4�E��q�w| ɘ��V}pkY�>��7�����l�N�=������K��e�J���HG#S�ӭ.�ʡ� �-�V���@��-�P�чa��!�|�o��QS��f(�XeD��.��Ia�Ő��#ά7W��d�L����kOÁڰ���d��m��؃�z��_�6�/L�D(�i�׬�p���Լ�,"���}�V���f��7勍1�n�ڣV�V�����2�t�6�㩱n?�0�$�p
����؂1<�7�цٷ|��R���o�-�.��flL<�5 ez'��-�#��ڝ����;��ޠ�b��[`Ae��ufߓ��L=�X�� G׶0�{�����.>��i~�F����;T�E�a9�a���-���R��#�x�z��NM��a�ާk�SO��Lp�N/V��4=`����RJ�.�v�{sɖ��3l�r�H�澚uA0���'_���(��}���ON�r ��V� Ha�~� H�|��G!y�z�\��x�OIz&��F�Jt�:�6���SQ���FA�hD�E(-Z$�"���0dNI:���z�p�w�x�Emo"CG��A�F�.�� ��������jң�� �/���WHcSvw���� t��ۊ�Ĩiq��:�]�p/;�}HA�L�5Cs���;s���/����Kxzl{�>�gp�쭯M&�.Q�Jg �[
�z��i�����]��`�b�1��.݅=)��S���+\ր\�<��/4N|g�\9��:�E��7�9�a%��=��e�T3�_��>1~��b��T���h|iZA�U�%h
�;з�M����^���}r��"�z�%>���h�Ɩet��c�Xf���;��c9}�.�6�
���
Q�5��9��9Kx<���!;��'W\}b�T$���5C�D �q%�|�����X��+�*|>T�]ȯ3?r���Yے O���-�n$�R�Gd�Y�w�~SEv�&��S�������KkJ>��ɀ}�㖱�
�!�#+���L�U,�L/�ru����L�c�H���~�,����mG���֌�eIt��Ԍ+��8�B
���"=�xTI����pi-����"�����V�F۬7�p�f����Z�c��Nd�R�c�c%.&j>��h\���� 9�y�p�G~\sȜN���'�;�"f\)>nI����C9���/���*6�8�O=��]q=G��y貏�xV�B��$��kc�91O,���(jb���#��潎
,*�ߎ]x)T����YBZ=ߝ���ఠ�<K�ۧL�22=ˁe����!*�x=�,|�y8�Z�
!j��
�TaaL�|.��F�	!G���P�[�2�!�T� ��w��7���K�����{V#i�ol��m��Ew `Fy�P�ٴ�����n~ ������;�{�t��_u?).�u�@��r�@�����L�ۦ�I������n���%�<�wI�E���ޒ��c@�.��	���v��[b�<�yu�e�:�X������!�(:�~	w���(�j������!c� ��a���8}��r�cu��=��~��y����4q�	���hQ�A&�3�1���C�o1����B��e�t[��Q!�R�i�S��Y�ʝt�|h����������9���cߓ��y�v�=���HN��i6���OQqr���g�	�ڍ�LfJ{���yߤ�)} ��u���f�
>m�鹰�އEf2���U�-�ΧHĿ��{��p�<}���ɩG"H.��@d��VB���Rm�J�d���y��ƃF�F�o=��VJ�����|�� ������d�nU��P�v��%V8�$�w�&:������8FĠ���fz0�i:4J�}�P�z���)�!|~teE�K:������εD��-���8�D1"S,ڀ!��WN=f٫�@����b����^b���	d�H#��3Mw�a�H0�x�h �x�z�