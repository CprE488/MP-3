XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����;�z؉&���z���)M��Z�bŘe���:Q�����]����y縉O�t��֡Qu���1�g4�Dv`¤|�Տ�o��:� ��h�%���Hڰ-F��m_{�jtm����N%��?����3�� fc9AYǗ�M���n��^q8s����6F�o�NADŐ��l��D�!~�m�o;���=�K5�6}V]u���P:�|{��fj~�c\B���n�w��霌�,�Nm7U$��4�J�d	�o�)�g��JV�%���9�_��\.�D���/�G���K���v�;hy���,4���z�z��]fK�ll�*]���_�q*ib�H�,��=���o��E�f��S�U�����\�⽊�9��+?�7gXQ���;4�>��2�ۥ`�j�N����a��Թ �}�O]�+��m�i]AQ���CEL7	���Oh�l�/�6��qL���\Nf��b�_�=�"��oL��=̓�C!LED��xq_>�5.	��z�<إ�9�'�B!�i�3K'�:�����r*�:��M�d,�V�.��᷎��{�M_3��Ty��(�֘��+��_��4?}�)�V'/���w9ֹq^A �MK��Ԋ"��Yşk|7�=�b��5�L�>q�9�U:P<��3$��X�w�=��i��!��Q`K�� pҷo>o4����DQ�F����3\cs�k�y�G��_x�H� *(�z4�u�}�y3JFX���Ө��9 =E4�(+�_>aH[ۿ{�PXlxVHYEB    5fea    1830��/"Jx��Z�C�vko����|���K�P��m	�S%�TY��L��>�٠\~�b��W�Fٙ���Tp�b׺D.�N�8��3c��ʫ�	2e��#�x����8�����
f����BTW0��SAB��e�cD��e�8�k��!|�����ֆ� 3ii��I3��CW�	�IPY��5��եM��e�\*��|��>Q!Ƈ'�e��l�:�O���k���om3��w�Q�f�=� 2ҵ�9�|׵P�cLe�1��e�:K7�'KFF�l������P�6tkGj���$����N�����M��Djhe�f	�H����v�5��N�����9�����iftҞE~��?и�PI�ft��O�׺19��OGE�\���ࢥ����fX���=>�W���H���"��n�q�yо�aVF�Sg���/��B�0�N��q1��U�b,����Q����'垎�p@}���1<N6o�����@�4l� ����oDU<��gj�N�����
q��M����B(g��Sz��l�݌��qt5�Vi��<au��t�f���̨�$ҤZ�)^�U�������9��EcG�o!�?n��z��^����Bx�<��ňB}�IwIUn��UvPer�Ծ��c�Z�
h	C�úf=�W��s2��_no�7�0��⁣�T;��p �?ä�c�&���ߔ62Y�z��D������`�b5WHwP��:JD+%jA$�Ù�pqj��F���L����Qn,����R��r�>���SQ2��%M�>%i��~Ӹ�?�K���n��q3aV�r�x����	`�8�X;�������p"Ajδߜ6Q�N����A��ː�8�E�G���G���]�����pN����!��"4!��a�S��M���K�@5>J/�w�4{��i�&��� ���l]���D������4�2|V�������55�������@���ѷ�*�t��B����S@&��J��% ]-�Y�Di����L��p}'7�Ɇ�RO�$��e2�43Z���U9%��=.��^��`��?�� �r=���s�a�;��	�T�e���Y�P���J�;�"(�� �ߕJ0��S�Õ[�f�O�3�-��c\����y��v��sP�&���lKp�:FC���9|rȘ�
�����Dw�V�����-"8=3��%�a�x|�^���6p���h�o�w!9����_:SW͎�.�F�w�D{�w;M5��n#m���2��� ��s'��e3=��p㔛�ƺ��ǹFNC��*�ռ.��嵝�2{CFk$W�1�^�p�G"!/�\>�Om$�����ȼ �����0q���?eUDoB3����2=Ώ-�d�O�h��W�w5������Dm)trY�W@;%����'���+6v��ӓq�sr}�Dtȣ�j���'A������� P6�*�"��;���#���Τ�O8��- p��� �n,Rk�®��K��v�Mv�EǑ&s���`����O"��,9�0�BY��!��t>��8�$��JP��N��G��������sY�ҟ`���-�M�X�*V�x�Ps�OJ_��x�٘u�,��x�������M��;��rpI�|�H��K�(J�P�nwF�m�_ �Z쬖�b�O�0)��v��bI9u��>k�d��WPn�Il	��ԼC�<�W$!d���Q9��RO2�iP�1XB����?�MbV:x�Q��jwa]"ogw���5�$���߲L� �@�K��-��p�6)�P�R��Β�d@����)��̶�Ń�*v��-����W��G;4��s!�$��l{1q��}�F��Ԯ� ,h�!����rϫ0�fk2�#B��hֿ5q�Yf֒YF�i���ڧ�������?2��3�;u=�����:��7S8)�O��M�CdI��kT�M4�h�}f���Gɏ�|M��#��#8p]cC�S�mswɴ7T�p����;n=sƕ?�Y����5Z��S���`��2�pNEA����\68�� [F.�P��붶���->MC�BC"�����T��-����#}pP��VҰ����|B�����֌��T��9�wkGN$d��ve�\)a����6����F?�nF�I�D�Ԫ&��9�c5���
z
i�	�7�8���沈��}�	\%4�# |8����v���?�"f�N(�ټ��?c�B	�tloH��jZ� �_U���m�Yn�o<jhݚ��C�Yg��P��A����X��^�9@DN�t�1(+q�@z'o�R�C�쮋�I�|����^pN<z��\� � 8�R��XG&r�e���*��sT�r�7~�5�i�8Q���S�Q�rY�N�g�/�LE֮��lؘ�p�+� SDk��#i@(e#�q	/.s��}N�$���PԼ3��|�խ5��5��W����l��b9�R��Kn�O�k�t�_�^�%S���{�-zm@�fB66��Ҏl�ތ%GUh��^U�h��Q:�J١l�꘴NC�aا'nJ����`y��UJE�5�#�%��˥?���a]M�mj� �����;�ξv�����`���#�0�gAg~�WA��0��q�ҋ��8��آ������p�#0����⅔�͛��ér&�e����)K*U8�Fsf�+8G�Q��Ujև�1C2�=�H�I��N�:��N���M�����0'���4��.f��{?�����~�$�%��@��!�ԐqѠ���oɦB$xw�f��i2�q[?+�lͲ[�`���!mH\����/���l��mJ��eG�9��9'w�
��	���٧4w[���{�C9D]��i@�PX��C����t�`=+䙕�j>"	'�$@��>����
��.��}l4��{K��� }�l���Mz���_�%:�=��K���<娻R�)ˋ�%(�^�^�{AH�A/u��g������H��=oS&ytWeP���%*V�F��>HYs�qU�}��h��]6?ŲI{�P���%�k�4��3��FANFN!,�V|����X'�Г�y͔��h0]��|��[GZ|�kL���S�n��1�{�� ��%�52_�x������NW�&q# ��*K� �H���ڿ>��L�����.�j�������r�zόּͥc�0���aTZ��_�k �D��`��E�Er���Lՙ�4Ɣ�����vy���f�W"u��Y���4���U�!����F��d�&(���g�k���[���z�J�/�`h��jD�u*��_�?��_�d�~fr8_pW�b%�4]�"?c�ia%�M�=�����w�d7+�tr1�3��o��'���A�A� �|�5#������c�iK�PWϤ�%��R��_��C��6H��V�g�e�$�\`3F�Z��v�j��#?�J�� >��5�b���3ً~��@����{ز�����/<H�')x���-q�E`�} �@>h_�eY$����2��4m�W���( T��ӑ3kU��7���Ng�w�f�^k���쾮�dn��6:+� b���_f��V�x6Qܝ@Qm�iڸ�o|��a{���T�s�w'���+��(FQ��@��3�����s?����OI�/����� m�m7�Z<�]U��5i�N����<N�-�i���[<�t�	}ŷ{X���BF�(��i4S��Wt�Ua&����Ios��fx͗�8T�������5S>��Q��k@�CY�؃"zm�I>6Ŷ#�tn�̠t���z2%<F����A��Et���8j���K&�����PC���K�Q�Vר������ 9�L~�Б��By�rB���W���S:A|\�F�3�W]Hg<��i�&ch�R�l� Q����[kv��5�n6�:��z��Tw�I��C��b�:��U�g��b�e �/�I�\�� �s%��d�>����[蘗�/���(��
����d��6��LD�v\�q���hO��u=�)	�ﮧ�홨��(#AKw6*'m��~iMg�٧�љ$���{�_ʈlL�#3�=�%ۢ��)?�C�4$���ѵP@5l|�y�ZU�����V���]e�bw�KM��D��fvs��b��/�7�>u숀
������Q���)=��e�L?k`2�L��!vն����Z���e�+�S$;��ܑ��㚓wk�'�ϵ�ס�H��	{8q��������Vf���ۧQ���o�"��מ�H�z�x�_S_�^����nX~���/�*�1�Y�"\,{D.b��l�!�T�]
XG�"[�!��K�@ZW��I�0 �?X�H�}[�o�}��W/p�6𢔾� N��^�6��������'�����|���H�HO*z;�7�զػ%|��#\@���)iX�c�̗����`+Y��H�ے��w�~$)��!�������`i�=�m���KƩY������o�8P�1����Y�w�M�v!���L�~B�������K�]�	�+��+yD����K���
d���
�Z�ϰ� [��nv7e�ic��K:a����^�2�P���{�<�8� ,��%喻M�jۧ��ﻟJH�ڡ����-t�kt1�ù��<��"�`ϖ-�C|oI�D4c/N�w��Nz�lB�p������U�饨udjJ��O��=�o!?�+��^�0l�fz���Ǫn����K<,���)�LG�E�w�FG�'�R�3SG6D�h���xdǋ���z۳մ�Z {V1� �梍�]vo�}���;��l9�V6�+dW?
S��1"xN��]��m�B���S7$��5j������0�M���w0jo�/��c��~�*s�W�ԒJ�/*���r�{%+q�q���2����1��O�v�^xq�)����ū�fD��=�|�͡>-M2Ks�t�Vm��Ә�|� ��?��൳��۔<h:��m��a"��ڵT4Rq}:z����)�Ls�� R��I4���jI���B fx`�gjX+�Ļx1B/���\��a�wXe�����{��85f��(����<rL �o��E�\�g�l������Hd�=�HW��ؽL?3�+��5e��!T��/�P��ei�ڠ���\�Y�Y�C7�)�|T� 'R�a�0A��'��Q���Y�T�d��}`)o|i˚%@���o�'�5}��}��������/�=�.�%-�K��L���Ջ
G7У�*��C��"ڴ��z�,�[x��Z��)���ۧ�<Awq��&�Sw𢦩*(�|*�3qF݈�w��!��ǫiӎ�� �N���2BR�`~��w�#��H�y��L8�4���{��~dڀ�3����|`�	��&�$դZt:|�ۏ��LJ�jXi�3Kc�,�:z8�/4�fZ�����"�zK�d(���(���S�J6n<s�s^;�|;dF����ۣ%^!ՑŌ���OJM16����v,#�`{=���I~����f��xc���)��'r�\��f����n��ҧ-c�g�Hܵh��A1���Ƨ��F$m:|i��[ӗTB�ul�qLזT���Td���ez�%M� ���M<�O��_=��Bb�&�@]��Z{vV��^m,p9�Fs�~l�x��E�"�|����� �Ȗ�\˫x?H�wQ� ,��)��u̞3z�f"�: G����|�wR}�#�&�'r����ش�+�s�%V��r���e�%����k+���n�U�M'��?�.psY»��=���r��)�*	!�*[ds�Q�՟��A!�d A�Ǿ����>�߹�����$N�,)�(�B�\����n�1�j3d�ɢ�����;(�׽	95�?5
j3�%N`l��x���4x	������� �CԀ��S���K�����3�0�Q�p��m���H��d�D$�B��6��'Czl�z��W�˦�S��l��g��P�@~�{�w�Qd�-|��s�����!�';y�i��/|b����}9
�_ ���`�M�T̨�vt���`�yܿ�K+V