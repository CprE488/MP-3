XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������&�o�� �R� �\#�c9L��8�AH��G�Ө ᥷�l���D�&_�+�K75���}ky!��K�D�X����;S�K�W�h��E�j��@�b������T�d%oʧ?w"�n�����[�)L�	R�~��t��Y�<��m�������A�P�v9�J��%�z�����P�=W�����V��O@�ז�oZ�^\����1 0���Ldqu=kJEB 	��$en�[5�<#��}�����Q���f\5/�?�} |H�6��ys̫�R_�B/���d5��հ�BפL^�U4�^J�6|���E��}],؄��I�،�V�yͽ���S���r�KecU=�W�d�o��^.G�u��R:kXZi_�/Y�V�!=N ��/R�wL:Ћ�MĻ���q�EP|@9��E�Mx�Y_�R��yRW�+w����p��d�����$�_fUl��΄�.:+��)����IZ�hz� /Om�Y���%���B��S�M�`b�1��Kf.ot7D2��Q��U%�RS�V��T�q�X�<ƫ��GJ�)��p��+�
������g�P�3��N������(�~n������7�3%pT.�j���Tǁ�,W�<�8�	�6�U��Ӣɜ���v���+I6��ֈ���ޢ�}��7�`�+	��D8P,��}y7����Ԙ��9�A������
��B;�P�	r��G��4]�sD��V�V��8����
c��~�sT�<6U��n�8����P�O_;�5�XlxVHYEB    5e2b    1530C0��E���yi*mƍC�bDNu2�L�3����5�O��=�N�Y�@����:��v3��	�X�+� j�"�m�Ip&F?�g!%� �z.,���^?S��'��oj���,� ����S�����Pݖyӏ�0�Y�O��G�[dD��dE�aNx�FM�="/&Jl)y�H�$��A 2`|�)���S�pf�½W~��jo�q��k�@L�>lP�R�rh&1�r���"hV*@<bF��q����9�n�;����4O�v�`�'��5Y�CKuv0���a�e/���B\�aEZP#[�^�֏��3N�hi��Nu\Ɵ�y�g;`��2Z#���~N�!�j@�W�ݼ�9.� l�ѠI>a��|��5J?'����8�ՙ�rt�p�#�2&��/!��'�S�ߞGd��x�� ����<�������sP�ρ���]�N�n��?�o�C��r��I�h�[Y���V����O��k�X�� �H�T�&Pw�*�A� ����FOߤq8�[�phF�vb�~����Y[=��5NI;�~��R�?5��x�sh�!^Y'0�k�����ǂ��4�U��� ��n��sU��o���]4}!����ַڙ���o�9�݌<c���8J!4���.Ͽ-��8��"�B��m_,K��D�kT��y#x��ǟʏ��۞?�I<�&��nO�A��~��H��⇡��LI�܌�Hr�֨�?���3�C$�B*����l�Az�ᰥ�h�P���װxH4w�/p.3�Ѻ�<�$Ց��j'm�QIo08�/u���:��%�2#�p�#�UY5���@��>S���Kar5*Co"��8�G�B��[�q�%�V&�&+�x#cOG���69L��&��"=�RG`��6�]>���Ō�wC�=/�ũ(�סT������ 8�t7<j��D��3l/�#� ��[�4.V��WU,n�����l[M'���`�-�7}�Pi`?Y�%�YB"A�`с�͞�P��Hi^`e�wZ����G{�HR+8;��>w��[��� �/C�o�c@H���a�egᤩ���C�\z��y K 29y~�Y�J,',��ui�����?�����1��/�	��;;����� @�u��:�%#c	^��m��}1OR��U�֡��Ò��$�����b��T�~�23�V�1�{j�J��;��E�GSf#�a�F�w�̻4�i��h(��'^����5�	;1�X0�����2.�ySh�z���2�Q6�A�5/�Yen� ��F��(qF]����+��.%m7��UQ*i��_�n��P�^<mIr�FMf5��7�u��i[y� ^��?���#�V�)�,��3l��C�Z��,hF, ���=޺��7f)S/]�ux�B�y������wVZ�?D�0�UPj�"'�.c��	��k��?pg�R��m2�
0O���J:� 'b�k��X���z��)ǗQU܏��+zQ&O�[x�$7u��nwtʒ��=x���#:��׊*�XҊM�ْ6d��?p>$�;ƿ��g�1eH�OӘ�a.w���b��)�zX���!�2 ��o������1:)+��d�?l@��kh&F�%�ۻ��ζ���v��l�'�ʛ��<���Ν�=܇ʴ�;\uWT���H
C���%8�c���{�L/�+
�C[� �+�T��QrV�ůLU4�E�O��-c�1���׸زC�A������(��"!���R0�L��=奍,����	&� 41g=��OQx��$�	���lN����s���_��lʛi���~b3Ѫ�h�4�A}nۖ�6S�o���yE�(D?������Z� r*"�Q�ZvnB���WM�n�
#�u]��(�����i,�Gh�Yk��H)$�Β�����A���D����may�y�s�-�.@�bX{��R�"��b�l����ob�p�'�8�4Ԛꨉ��ǊJ�6����-ƅ.KQ��09�`R#R��Hز� w}k� �l�b�a3a0�O��U� �0U�o���K���o����ܫֳp��A�c�7@����q|`v���M͔���Q}�y9�I��kW)dL�2O�u;��QkY�o��b�A*�=C 0*�'�p�6<�GaR�z@eR2��_6�|n��(_CS�'}�9Di�g��הC�̃^Yc��������ǯ^T�
P�9@��5�H���f���"ۥE�뜌'���ͨ�T�1o�]~��:�$�B`�D'&�hC0�E
=⛬c�����X�c�?S�E�S�-+�5͒����))$��P;��������!����/���b�.@�Ƃ�M.F4~�	���N4�;4�~�=MG�K�C��&�
"��JT����E5����cT����B �M[�Zt��;�آV,A#W�f��>1��F���Hx޻BT�8�Y�(�Sxm�����R,Hc	�����n龜�z�Тt���*Y��93�5S�89"Σ��t��}�5Q�,2���F���G�6o���]��0�̲�?�K�ÆD����5;�:�ܿ=�[� �uY�_)�13���Z!XX���&�m|euTY4㤪΄�
�`j�d�er�h�ø�S�z�.+�¾�f:�Iu���.n�Z�V8}�>!s�oY���Ӽ_�H����ѲŒYbw�Qj7��)7��x9���m��e�#��6�\���c�S_`!d|Y�{��H�����0cS����\�^f��I�_Yӷ�hK���C&����2^a�&ցF��|���s-���kb|���Ty.6�U���H3O��g���/w��?v��ӷEF-��F[-@��h_���^�rv��t<�jZa�b���p������@V��}��e7���� ��(A�}Z�����N�����h��qZ⋲z�G!a�~Lň�r�x|�{*$0=_}��[��b�������F��ԉ��=���|e�D��KP��h����:]����4<��o3���+�.�x֡xq�ᅽ���֒�xG����x>T�ה�4��V1F�A����0S���w~�����r���m.����Aw)�c�ͤ7�����e���ԓˇ�⩶��6�	D��2\���g��]BiRpJ+[d%0�=�����r<��z������\��&-�s-�p���h�b]�y��=�a��	�b�E�N�]�*�&ehx�y�p8��� ��K;�(P���=�7=�q`]5���M7S�x!HAq�~�Ⱥn�^`����J<涄C���q)�S�	o��KZ{�6��ƣ��۷%�E5<�:��C�5`q�a%j<�==<���]uQ�e�pW�d�j>�����PĪ���m�;�O� &�����	Yrt�c��/����S�{c5*����U�px7*�h+&*��{��IY��	9���fN:�-��B�)NZ��� ތ�f=�e�B�i�ۄ�J����VV���ޓ����)�9��v�C���p$����yW�d�:��% ��!̚�2���3�G21�谆�7��RH�L���
�8vnF�қa�|!���D!|L�eK����i�+�[�Y��.eA^wo�~�=��4�u�WsT��Ml���}�X�����|>#��<,;��l9�+�*	�I�yt5vV�NKmʥ^vY��6�vmp�^�OL"���km�����>�*����d�h�!0�r��6=�W�ș�k\"��7!�"М���3pQ�L�M��W�>�~�Y��w�Î��.�&۠a�D� &���8	O��&4�KT(�*�� ��ħT���>�>��Z��eE��)~q�����u�a�ͻ�h3�>T��� ���8��D� ���<�U����7IW�����V�^!"�@mh������!/�/{g��v� Y�'�ô�{��U�Vm�0�-�"@�����][C��`^U�7�Ȭ�˺��Qqe�Tɱ�?ָ�=�;p���4�������ޯnԱ��3�W�o���`{��c ��p>��2
5��*�ϠQ�쯘����h=�#_�ѐ��35�h�>$�;�)G,+��:ڥU�DM�i,8��:�x�^��eS�fL���͋�`A��Z��@G��-�BK���_�˥��!�N�������}���6�Ś��3�DA�"�� ���f��E�����p�Yu�5sT��4�KOO��c���a�?���p���Џd��P�"(υ�D!��U����L�p���� �EUGC-L�5����~~��%kk&D���v=z���)�X���y������==yԌ�Tp�x�G-�{��s&��ް��j"�p��V�G�C'X["����P���7;͕WU~�iuS�;�k�~ڱ ���F��tgq�I�N��Z�e�WL��/Iv_*�w��o/��v�q��x��J��D�g<���<Q)&��Q��O=�U~�p��[L;���&��*��rc�B��k���Ή���7�����$������0����H�SU]I��.B���ssdMP�����A�&�Gf*��1�����[u}$�T������C�R�ڴ��=*�h�=�/��N񼞨s��r�+=*���U�ï��cy�d��#F!`˻x�5$�H�L�w󼦯cr?�n�v�Nym��t=;�A�[�׉i���>
Wj��i�>��7Z��g|�W!J���ð���U+&8e�� �H'F)
P������uoC��O��fU	F����a�h\��4��kw��Z��s*�ņ}�1_-IY�dp��v���BÜ门����w�`l�&�8m�&��]�M�EЦ�9l�8I�N�� �n�:(c��!L�Z7�!��L[>���C�zj��mK�"y9�&!��B��i������1�`��S~Θ�u�#<���Z��b7���?��b��o��)=	�-��>k#�[�ȓ������	1�k��e�!��>��S����S�h��i��9���)C���͗r�Q��1∥X�l�IF���NF��?�������U�
��`�ő�����Y����ECHʥhvFi8b8]* u'�m|OC���q}�"硾�0�,&t�
��J�1��@MwDC�%�©��0���&��:,2����\��7����m�<��j�T�t�.�sr�\��B��<��~�[wU��<�5��)+�����HŖ Ne�EDB�䫝�~�B�.�烙-�m4g/�R#���fg���f⢻�O%s�[� �(�_[i_��h��?��F�镞+�z��#
LS���[x:�XA�8�X4$��@s�I����5���S��V��,�|7�