XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����N������o�R�>���M ����Q1�O��,�Ө�(=��Q��O�eE?+˝�`�|��f0j�i͘MU$�k��܉�}�]���U"=��˧�_X�?�IԨܲ����߱�E��������Y�c���S)m�U��lOi�L��R����	�{Q�� �,��տg%�e��-w�8�=�o����O��.�*7�P�GQ�_�ט<��7��,�,0h��ݓ�:r����]�	uK���Ҙն���v$G�*�'a<���U�JRAxQ�r�h�%�������P��븿���
qG$X�I�>~M��an>ՠЕ▫�
�� �ͷ���F�=��NL������79�.#ew�}�X���ý-��"��T�%)������	��L���1��7��;i�z��xPm@�����D��PpY�)F+2�p��
�4՗X+r��Z3V������e��w6�d��Aޅ�ʖ�"e���\��
e��*�*�q�衶Ŕ���mbx?�k�j��z�Z�K>CfH���.i۬H�F}�x����\��#��u�f7�� �!�g�_��͋�W(�U8�8�J��3?��RiG�D�����S6K��X)u�fw�����Ϭ,F��?�I�žq����֑þqɌL��<��_h���N��̓}�\��nO �+�9�o�tz{n�� ��DBs���G㩙��d��J2�§�ʝ�]��r�oJ�Dk%�L��+��,˝6�*'��dgf��#XlxVHYEB    893b    1e30��
��v��Xu1 �I�ujWy��Dk�>$�Y�
Kd��a�и�u]d��
��T�dY��J��[��]Z�z��b�i7�:�����9Hb�#�`���6���J�	vL��{/i����sngy��_|hh|�����Q~k��N�����\2W׈�a�찆�3h����+�> K�kӥ�/'���~�XE��z�`=b��Ni�R(�Q���Wo�|S�Di[%�?�?��O�K���%Qg�i�NԪha,�S8v��������D�W��3E�3Y��޼�py���
�����_�K������
m�Hy}?�g�@�A"M�:ӱ�TጶdN�_;x8l�-��U���f0�oo��� R�"��E�>��{rm�p�G�{~��RSՒ���H�~j��2
�S�$����j�$Խ�2���<�b3�h��(>;RW)�FU�a��΃E�~u�iYFK[CL�noL��D�{L���nR��&ܻ���Z��7�ffžfy:����h�~%k�{�T�)�ʽz��)�r>bz�<Vkm�eN����Pimo��u�{ǆ�C
���$�����a��0�F�CZX���;�����Ceu+�j$:�Hع�]e�*�ے	&"�^��E'��lN�"?As`��ُ[l��-��2H�\��z�43�0<D��.�0�nQqiw�(W�<�ς��G�J�qx�Z?������^h�-�p��0�t�
l�@ٟ��9�F8��Nn���Ve�Gh������U)3VPf(̞G�IEaY�?��N����0R�@. �t)�>3��0"����	�W�:���6㳭b���f3�[�.3PȂ:N�ڣ�.��*��F���%��/z��xx�G#��4:؛m�{�I��bش�Ԡ�efJ�"�k.]*VL�C�s[ �6�j|F���,��u
����t��8����p�(f%���T����Y�N�Q�k>�Ɲ��j����t������@�,�&|g�H}��{�x�DT�Ό�w���m�S,/������l.���:�z��dc�]��\�����m����c��j�KX�����<�*q��Vb�l�vF�>m��!W��
I
�� � ���ZW�QI-��߽>��x<H`�#�"P3\��ˠ�o#i�Jwˑ�	q�H�U��խ�]ay6���d����7�IdGx��:��"�'Ԩ�\��P����Lg��W`����ۍ����mι?~�+s������D���Xj3� X�;ֲ6t�C�ŗ؝�pY�(Iz�����O�s�;`�`��\�^�/����6͈<��V���P���*�4�@Ѯ�Иh�ͿO=����T;mɾ�S��4�%�A�pcm��B0r |���%���v���2$��/�V��:�L}�R��\�U�U>I�/>�ٱ�o�����V�E^(�8�=���*&����g~�.Gd+I����Tz�=��֥J$ϽԆ�%0Rd>�m�T�G(��U��~�Lg�0��f .q(��k������1���h�26���3:,��Rk��{���Yo�����.���1-
"(�y�;�S��aqG��+�e�k?9�6���(C#�e�Ֆ/�Pl�����Q��g��<� �2p�WHi��g`ZK��$�������!����	�Q��S r�.AhL�ڽ-tX<����:�U�Ǘ�y�#d��n\+gǅVQ%Xр�{!j��'k~T���~|t��Y�X���'�F'
Qs�l�Kf�.�����A�N1��N}���e��xBl!H�ɗo��R�K�8Tn5��	��ULR�ތDkh�I�����%��z��4N
x�_�u�S��g]w��ٰ���r��1m�s��Һ��)��e�}b�L��l��9�oe�4h@�ɼ7�|
Q�A��=Pf(�T^;���qlJl4�?�U�F�i�WX4�D���
���аh CzU+jm�`o�����ZEw�!܃��u�Z��W�68Q2x��
���?%F�~�L�R��֞Z)3Јl/[4$�6&��y'�fVO}�]�6����Tq0?�<��b�x�>�>�.�9]�A��\�G�f���p2D]���H�EY9��:���+�����/��UZ�h���ء������D8("ˑ谳���Y�z���L3��w�ʈ|��AB�������;�f�<�q$t�TX�l�z��,A��`�Se�R06g��0�VR�g��0�Sq�q��ᐃ֕�Nh�c�tW
����ԭ`�����ܨ�Wx�u�lv,�@�7�lݼ{���Jn���C���J�C��X"�L��p��r$�GmLz�2-X%�
�F�ț�u�����V����rǺSE#��M3|CX���i啬l��D7Q�lϡ! ��4��@����t�y9���[x&&��1��Ƃ����6���̰��r�zC��㨢>��>�c¤���[�ߛ6�E$/��}�[�+7�v'��Ѧ����ǗL�k_��������f����"�,݋6�"�E�ˈUz�l��ov�Sz������@���q�� �xR�0ڳD��VZ�nE�+���k`{�
��r�e�Rq�R��)�G$��j?���8a#����c1?6Э|��E�}9^��1aAɣ���%a~�q��XG6l�_ˎ<�O�,��?&��p�����]s��7�c�CR��i���FW}!51e`��Ϊu�/�#�(f�l��b���T�T]>4tiU�Ͽ����ܼ?�Rn���)�'��b2.Og`�ly�!�y�����+��F�8*����A� �k�Q��졻��o���0�>����k{����ȷ�qË:C�	*���tنG�Ý�c�,�7��-����S�()s뱃-䵟�Q�R���
�0�>Po�!�-������; �lx�١*t�f���1F���le�Qy:TE������7a ��#�!/By	Q#M�t�g�sA�$�}���h��S��R�_�Fc�JM��vv��|�ٜG/��w���_̃�Ǻ�����fLF�k,S|��R?� �%Y����L�����T��Eg�'!Ond��M�����pP���F����(A?�*��蕱�M�G�R.��5��m��k['bjZ��@{�_1��ܢe�`�`8j��sI��1�IK4m���m�L.�G�8��z��R�����bٰ�쐈C�+�P�+�����c��E�n�uw�=����킣�-dZ�����>]�5?_,@�Q���6�a�Z%��D;V���,�*+���R����+��FM�u!0�N۴���螶��,OC#M�h����L�j#�������%MT�m1��Sw�uK���R��9�jR��aB�@U%'�¼{�!��ԦX}�j]󑍽Xv �mg���#�^���4[Y��+��:�;���m�_ke�Z	K+s�bğ�6K�߄�X��*�S�O@�Yi���)P_W=j���DQ�g������k'LHH�!��L$ñi�0�<
ы_=�>�l��GHH}RO��ɡ4�~���R�9"�5ur)2�m5�G�N��©��k�Ķc(�ל�d�"���%�V����a��,9ح_��\��w�'�v�΃{��]�"f�t]7:�1�:�_��[+�t�z�z�IC��Pfn]�S'1��ARfge��(!$�O��SH���~63�"1���҃��/�?�Ȼ5V2'G�J�� ��a�����)��F*�}����|{�;��x����E���x������f�e��y��@f��Y�<�/���^$�B�-,6Ss�j���U-�y4C܃��lU��$2����VPr��B���:�4Ȉx�ї�H� t��ZĘN��
`�c{@ ��o�i�˩�@���os��bxӢV�1ڜԏƱ �iXN.\���UUZ�
yS}FFa뮌ulc����A�w�ճ!�b
�h���3�(:j� Ф_틌&�zK�DrR�|�t��Yʟ�?ӻ��҄���f���2�g8�r"�K߱�u����	���Z��zϿ��u����mY�A�L�q$學�jM�a��}�4|����ױ�X!�X����9R��vC���+	�4���s�Ih�Z�=ul'�h$�B��Z��iM^����GV�^� '(�͆׽,g�RI�~ƈ���/�!���^L��.�	K���1�@������r�T2z!_�5Vci��T���1đs�昬�36�I5�cM�sL��V���?]���4 e�d8hX���mw����&��ӝ��9���<� ���� �N����`�	_{�[��^�ng�f ���Gx���%�^`�A@�O'�6" ��R�]J/l2b�R���z�	�K���vQ��R������8=�mf|h�zaim��{<�$��^��ي�P�..$2XS	�l�`7abWLt��(�[�ہ�+�G���d)z)�,�/�Sk�]��k�2>���3��=SZ�Fol���A�H��)���oY�ɦ��GŸ��i�i�{׵w�V>,!��J���[[4�V�#��bN�-_�7��縈@5�ڈ�vE/�)}����}������������㩸?AZ`(䊘ہ+�&={^d|�.�7�3-ʡ>i$r�Q
1�
Ft��wx[EZ�����Y�C?X^>�&
m^]���Z!��`.�]�(iX]�2��`<PQ�@6}o�*�@�᪠��i�2���a%��_Q`%��[��ݗ�*����M�i�r|D�";��|�^�� �k�R=�:�Td���(����^�L����6f������-�tQ��\ț�H�2���ɡ0��b;K������4O���Q<��q�����c����kn�|����ﱰ\��4�n�B�5��8�4h�C�vY��3 ��U��(Z5݌�*-΀�3�/<_�#��Ws7'�P�w�K��^ w(�@�ș�v�&VN� Bh�ӟ�@`Vd�4�u�M��՛��W
�������h�ZBc �RNU��͒����a�bF�	�¢yC�#���]���AX>��K�T�pG-Z/N�k�t���+�)SL�X�K7yXg�3�(���3�4n�رu9��p��f�X4w*�B���3�9��"�Ԡ�71�y�]�I3�R�gЖ�l,K��L��GL���-4=Eh����\�x}�,�OsmI�p�Ҹ8 L�]��C�� [=GeU$j��܄�FJ/��@�$��Y��iybЕm- f�P����F��.�^#�{�h�2
��Jl8P$FH����7pLL���P�b��ƹ<����(�JCrFlkN����]����;�Nt"�yր2���!s�!fJL-��tʝ�S��H*�r��Y�2j�����@�l}C��. �f������l3�O�~���+W���������A"QT����>Z^����$��_�\h���ƨ� ��:����qr|v 8���b��b[I�~rSi�9H�߄'��Q��|3Q�S��sw�yA�m��h������LH�9W�=R^�A���WQ�n�Qe�����/8�_`%�ʨ:�`}��x?�
���H�Ņ���]iJ]��Cy�\֟�W�ꘆ�&������DU�:G^y����q�ÉjL\�RQ�L�j�`	�ZRR�61d2���D����VIK����O�h���PsZ�*��l���4�^�:�1���ߌ�ahyu�nU���3��6�=A��ܥH��~�rJ�N4�Ǌ*��O˞��#�J�|5�I������0�q4�2��\J���SǸ	��V�0\�-7��5���>�����03}1��Jb�c�������0$
�9^�֪�v�֢(J����,{��0���b+�|�E1W����U>|S��F�j�Ň'w`�_�$Q7��2��B\��{��eIo��Ð�%>�'�
ޙ��z7�]��:�g�u�u�f3�<
���`u��%?�M���ӡ��i��I�SlQxp�?U���Kg7wӵ��N��#)i�cC��H������I�?�K��ˏ�ː���;jE''�bG:*VV�����alF��z�"�-9����Z�'$��.��O�)a�{�\�/~�~l������臂r�X�iK����{�iXJP2T���*�,Y����@��Ի18�՚[�d�O�/+ep��l�W4E'[��&0��i�_���ʥ�Gd{E�IO�A��ա��O��`�8�<�rj4�	8c������r�z�5xs��Nw�!��g�	d%$�)�ќ0�C�7t��:�
�Q��Lz<��y1顩|��Ȯ53�5N�qG�R������Ot�{��nT#Rüw�f���f/cS�[G��=W3�­b���Tf�>3��	<�[�+��(���[%$�S#�")�:�Aˣ4��;�9����|�
��h�}n#�f�з��(�G� ^hp])��$�"�N`���[��e\H�bU���6�Nň�"�s��D3[s0F����ķ�h��y�y��wGp��
��[x;?@LUH����ܦ��$�8�素����#M6nb�T@ښ�������whP���) ݿ�@���ƌHq�I�k��䫁!�šMd}+^���I^��,��=M��K�
q��I�adc,��rqF�DL��̿��i|r����6�̄��}ͿcW�\�x-�E���u��π�.>�1_;C�Le&��\[�Ux(�������W�8��2��U�gl��o>�΋qJ�u[���)����ڈߖþ恱-b�5TF�;��x�!�K_Ć�/��D�WJ�_�|(!����0=\�v���fQ��Nou�v�q|�� ZXM-ꈁ)�#|��H?qj���Ʀ����:���q���~J�Y��?g���%�wT�@T��ŵ ��\�K�wCo�pKG9��0qU:9��b�&d}��x�)0h��:���{�+�ۡ(`f5D�#����-�����h�ܨ�y�˻�R��E0�]�w�r|T��|��3S��������-OG�Z������\�į�97�攴I�M�o�Cj�zA}�nt�y��|l��4� ���fF.xPvTÅXH�D�����6İ(��B�f�%:���mf�1�՛���z͚�i<vu?g�/0'�~%|����_�Uʆ�x� �%�_6/M��n'6��%i�Σ�+�(6Tvq"�J�qB����T�5.��|�˕��#��kt�
�"�%Wz)e-Q�y��9Z��Rk�Z��R����~��Y�!%/\=�� �g����1����8�C�s��u�y�_W�$r ��
PgI�Uu� �>�m*��(�� #z8oއ��X�m�_(�����m63�!��S�1�1�/��cpB�Ni _�%�b��г�e��';53Lz�\��e�̫D'�����Hեp�|�C��y�,�1I����d�Ik����Q�?�N��N,��~���"�z�_rŌ���\�u/!8m��,d�9,�6cQ�x��+�;f*�_��XRS<�~��;X��ο�����5�+W�������t	��y�mg�~ /h�-Gw#h�`��D�|#���E'�m����S.<S�qi���m�������*�0�uL��=���M�w���T��SPg�>)�� ���ia��}���V����Mf��